module shared
