module executable
