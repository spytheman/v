module sharedlib

pub fn version() string { return '0.0.1' }

// Put here stuff that will be defined and loaded only in the live shared library.
