module live

