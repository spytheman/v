module shared

pub fn (r mut Reloads) load_so(soname) int {
	return 0
}
