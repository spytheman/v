module main

import zxyw

fn main(){
        i := func()
}
