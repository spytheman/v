/**********************************************************************
*
* BMP render module utility functions
*
* Copyright (c) 2021 Dario Deledda. All rights reserved.
* Use of this source code is governed by an MIT license
* that can be found in the LICENSE file.
*
* Note:
*
* TODO: 
* - manage text directions R to L
**********************************************************************/
import ttf
import os
import strings

const (
	font_path = os.resource_abs_path("Qarmic_sans_Abridged.ttf")
	create_data = false  // use true to generate binary data for this test file
)

fn save_raw_data_as_array(buf_bin []byte, file_name string) {
	mut buf := strings.new_builder(buf_bin.len * 5)
	for x in buf_bin {
		buf.write("0x${x:02x},")
	}
	os.write_file_array(file_name, buf.buf)
}

fn test_abc() {
	mut tf := ttf.TTF_File{}
	if create_data == true {
		tf.buf = os.read_bytes(font_path) or { panic(err) }
		println("TrueTypeFont file [$font_path] len: ${tf.buf.len}")
		save_raw_data_as_array(tf.buf, "test_ttf_Font_arr.bin")
	} else {
		tf.buf = font_bytes
	}
	tf.init()
	//println("Unit per EM: $tf.units_per_em")

	w  := 64
	h  := 32
	bp := 4
	sz := w * h* bp

	font_size  := 20
	device_dpi := 72
	scale      := f32(font_size * device_dpi) / f32(72 * tf.units_per_em)

	mut bmp := ttf.BitMap{
		tf       : &tf
		buf      : malloc(sz)
		buf_size : sz
		scale    : scale
		width    : w
		height   : h
	}

	y_base := int((tf.y_max - tf.y_min) * bmp.scale)
	bmp.clear()
	bmp.set_pos(0,y_base)
	bmp.init_filler()
	bmp.draw_text("Test Text")

	mut test_buf := get_raw_data(test_data)
	if create_data == true {
		bmp.save_as_ppm("test_ttf.ppm")
		bmp.save_raw_data("test_ttf.bin")
		test_buf = os.read_bytes("test_ttf.bin") or { panic(err) }
	}
	
	ram_buf := bmp.get_raw_bytes()
	assert ram_buf.len == test_buf.len 
	for i in 0..ram_buf.len {
		if test_buf[i] != ram_buf[i] {
			assert false
		}
	}
}

fn get_raw_data(data string) []byte{
	mut buf := []byte{}
	mut c := 0
	mut b := 0
	for ch in data {
		if ch >= `0` && ch <= `9` {
			b = b << 4
			b += int(ch - `0`)
			c++
		} else if ch >= `a` && ch <= `f` {
			b = b << 4
			b += int(ch - `a` + 10)
			c++
		}
		
		if c == 2 {
			buf << byte(b)
			b = 0
			c = 0
		}
	}
	return buf
}

const(
	test_data ="
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
00bf bfbf bfbf bfbf bfbf bfbf bf00 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
00bf bfbf bfbf bfbf bfbf bfbf bf00 0000
bfff ffff ffff ffff ffff ffff ffbf 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
bfff ffff ffff ffff ffff ffff ffbf 0000
00bf ffff ffbf ffff bfff ffff bf00 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
00bf ffff ffbf ffff bfff ffff bf00 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
bf00 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 00bf
ffbf 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 00bf
ffbf 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 bfbf
ffbf bfbf bf00 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0032 72bf
bfbf 0000 0000 bfbf bfbf 5400 00bf ffff
ffff ffff ffbf 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 0000 0032 72bf
0000 0000 00bf ffff bf00 0065 9999 ffff
ffff bf00 00bf ffff ffff ff7f 0000 bfff
bfff bfff bf00 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 0065 9999 6500
0000 0000 00bf ffff bf00 bfff ffff ffbf
ffff ffbf bfff bfff bfbf ffff bf00 bfff
bf00 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 bf72 3300 7fbf
0000 0000 00bf ffff bf7f 5fff ffbf 3f7f
8fbf ffbf ffbf 5500 0000 5fbf 0000 bfff
bf00 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf7f 5fff ffbf 3f7f
0000 0000 00bf ffff bfbf ffbf bfbf ffff
ffff ffbf ffff ff7f 0000 0000 0000 bfff
bf00 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff bfbf 00bf bfbf 8f5f
0000 0000 00bf ffff 7f5f ffff ffff ffff
ffff ffbf 5fbf ffff bfbf bfbf 0000 bfff
bf00 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff 7f5f 0000 0000 0000
0000 0000 00bf ffff bfff bfff ffbf ffff
ffff ffbf 0000 5fbf ffff ffff bf00 bfff
bf00 0000 0000 0000 0000 0000 0000 0000
0000 0000 00bf ffff bfff bfff ffbf ffff
0000 0000 00bf ffff bfff bf00 0000 0000
0000 0000 0000 0000 7f7f ffff bf00 bfff
bf00 0000 bf00 0000 0000 0000 0000 0000
0000 0000 00bf ffff bfff bf00 0000 0000
0000 0000 00bf ffff bfff bf00 0000 0000
0000 bf00 bf00 0000 0055 bfff ffbf bfff
ff7f 00bf ff5f 0000 0000 0000 0000 0000
0000 0000 00bf ffff bfff bf00 0000 0000
0000 0000 00bf ffff bfbf ffbf 0000 0055
7fbf ffbf ffbf 7f55 00bf ffff bf00 7f5f
ff7f 7f5f ffbf 0000 0000 0000 0000 0000
0000 0000 00bf ffff bfbf ffbf 0000 0055
0000 0000 00bf ffff bfbf ffff bfbf bfff
ffff bfbf ffff ffff ffff ffff bf00 00bf
ffff ffff ffbf 0000 0000 0000 0000 0000
0000 0000 00bf ffff bfbf 0000 bfbf bf7f
0000 0000 00bf ffff bf00 bfff ffff ffff
ffbf 0000 bfbf ffff ffff bfbf 0000 00bf
ffbf ffff bf00 0000 0000 0000 0000 0000
0000 0000 00bf ffff bf00 bf00 0000 3f7f
0000 0000 0000 5fbf 0000 00bf ffbf 8f5f
3f00 0000 0000 5fbf bf5f 0000 0000 0000
0000 bf5f 0000 0000 0000 0000 0000 0000
0000 0000 0000 5fbf 0000 00bf ffbf 8f5f
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
0000 0000 0000 0000 0000 0000 0000 0000
"

font_bytes = [
byte(0x00),0x01,0x00,0x00,0x00,0x0c,0x00,0x80,0x00,0x03,0x00,0x40,0x4f,0x53,0x2f,0x32,0x41,0x98,0xb7,0x90,0x00,0x00,0x01,0x48,0x00,0x00,0x00,0x56,0x63,0x6d,0x61,0x70,0x53,0x38,0xf9,0xae,0x00,0x00,0x03,0x60,0x00,0x00,0x02,0xa4,0x67,0x61,0x73,0x70,0xff,0xff,0x00,0x03,0x00,0x00,0x3e,0xf4,0x00,0x00,0x00,0x08,0x67,0x6c,0x79,0x66,0x95,0xf3,0xc8,0x23,0x00,0x00,0x06,0xe8,0x00,0x00,0x2f,0x6c,0x68,0x65,0x61,0x64,0xf1,0x64,0x88,0x06,0x00,0x00,0x00,0xcc,0x00,0x00,0x00,0x36,0x68,0x68,0x65,0x61,0x11,0x4c,0x06,0xc9,0x00,0x00,0x01,0x04,0x00,0x00,0x00,0x24,0x68,0x6d,0x74,0x78,0x03,0x08,0x1c,0x4d,0x00,0x00,0x01,0xa0,0x00,0x00,0x01,0xc0,0x6b,0x65,0x72,0x6e,0xe3,0x4a,0xe3,0x1a,0x00,0x00,0x36,0x54,0x00,0x00,0x02,0x22,0x6c,0x6f,0x63,0x61,0xa1,0xec,0x96,0x76,0x00,0x00,0x06,0x04,0x00,0x00,0x00,0xe2,0x6d,0x61,0x78,0x70,0x00,0x7b,0x00,0x9a,0x00,0x00,0x01,0x28,0x00,0x00,0x00,0x20,0x6e,0x61,0x6d,0x65,0x86,0x7c,0x31,0x7d,0x00,0x00,0x38,0x78,0x00,0x00,0x05,0x5e,0x70,0x6f,0x73,0x74,0x21,0x0a,0xb6,0x4f,0x00,0x00,0x3d,0xd8,0x00,0x00,0x01,0x1a,0x00,0x01,0x00,0x00,0x00,0x01,0x00,0x00,0x17,0x61,0x7a,0x59,0x5f,0x0f,0x3c,0xf5,0x00,0x0b,0x08,0x00,0x00,0x00,0x00,0x00,0xc4,0x10,0x0e,0x69,0x00,0x00,0x00,0x00,0xc6,0x1e,0x2e,0xbf,0xfe,0xb5,0xfd,0xbd,0x09,0x63,0x08,0x26,0x00,0x00,0x00,0x06,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x01,0x00,0x00,0x09,0x31,0xfd,0xbd,0x00,0x00,0x09,0x62,0xfe,0xb5,0xff,0x39,0x09,0x63,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x70,0x00,0x01,0x00,0x00,0x00,0x70,0x00,0x68,0x00,0x05,0x00,0x31,0x00,0x03,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x02,0x00,0x01,0x00,0x01,0x04,0x34,0x01,0x90,0x00,0x05,0x00,0x08,0x05,0x9a,0x05,0x33,0x00,0x00,0x01,0x1b,0x05,0x9a,0x05,0x33,0x00,0x00,0x03,0xd1,0x00,0x66,0x02,0x12,0x00,0x00,0x02,0x00,0x05,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x80,0x00,0x00,0xa7,0x50,0x00,0x00,0x4a,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x48,0x4c,0x20,0x20,0x00,0x40,0x00,0x20,0x22,0x19,0x07,0x47,0xfd,0xe7,0x00,0xcd,0x09,0x31,0x02,0x43,0x20,0x00,0x01,0x11,0x41,0x00,0x00,0x00,0x00,0x00,0x04,0x00,0x00,0x64,0x00,0x00,0x00,0x00,0x01,0xfc,0x00,0x00,0x03,0x7d,0x00,0x00,0x02,0xb1,0x00,0xce,0x02,0xd7,0x00,0x64,0x05,0x0a,0x00,0x41,0x04,0xf9,0x00,0x45,0x06,0xbd,0x00,0x20,0x07,0x03,0x00,0x92,0x01,0x89,0x00,0x64,0x02,0xaa,0x00,0x7d,0x02,0xaa,0x00,0x51,0x03,0x1d,0x00,0x4c,0x04,0xac,0x00,0xc0,0x02,0x39,0x00,0x9e,0x03,0x14,0x00,0x14,0x01,0xff,0x00,0x9e,0x03,0x3c,0xff,0xf7,0x04,0x73,0x00,0x0d,0x04,0x73,0x00,0xa9,0x04,0x73,0x00,0x28,0x04,0x73,0x00,0x20,0x04,0x73,0x00,0x00,0x04,0x73,0x00,0x35,0x04,0x73,0x00,0x0a,0x04,0x73,0x00,0x1a,0x04,0x73,0x00,0x11,0x04,0x73,0x00,0x21,0x01,0xff,0x00,0x9e,0x01,0xff,0x00,0x9e,0x04,0xac,0x00,0xc9,0x04,0xac,0x00,0xc0,0x04,0xac,0x00,0xc9,0x04,0x73,0x00,0xbc,0x06,0x44,0x00,0x40,0x06,0xa5,0x00,0x45,0x06,0x8f,0x00,0x57,0x06,0x12,0x00,0x3c,0x06,0x4a,0x00,0x34,0x05,0xbd,0x00,0x38,0x04,0xb2,0x00,0x35,0x07,0x0d,0x00,0x1e,0x06,0xde,0x00,0x1d,0x02,0xc6,0x00,0x33,0x06,0x92,0x00,0x51,0x06,0x61,0xff,0xf9,0x05,0xa0,0x00,0x43,0x09,0x26,0x00,0x3d,0x07,0x06,0x00,0x3d,0x07,0xa7,0x00,0x1a,0x06,0x50,0x00,0x3d,0x07,0x93,0x00,0x24,0x06,0x5c,0x00,0x27,0x06,0x28,0x00,0x2a,0x05,0x97,0x00,0x01,0x06,0x3f,0x00,0x16,0x06,0x4c,0x00,0x02,0x09,0x62,0x00,0x02,0x05,0x68,0x00,0x12,0x05,0xe9,0x00,0x21,0x05,0xce,0x00,0x31,0x03,0x20,0x00,0xaa,0x03,0x0b,0x00,0x0f,0x03,0x1a,0x00,0x50,0x04,0x2b,0x00,0x00,0x04,0x73,0xff,0xa6,0x02,0xaa,0x00,0x4a,0x05,0x02,0x00,0x3e,0x05,0x15,0x00,0x4b,0x04,0x49,0x00,0x39,0x05,0x35,0x00,0x34,0x04,0xc0,0x00,0x39,0x02,0x70,0xff,0xc6,0x05,0x02,0x00,0x27,0x04,0xc0,0x00,0x42,0x02,0x73,0x00,0x52,0x02,0x12,0xfe,0xb5,0x04,0x52,0x00,0x3e,0x02,0x3d,0x00,0x38,0x07,0x96,0x00,0x46,0x04,0xd4,0x00,0x46,0x05,0x51,0x00,0x2d,0x05,0x0a,0x00,0x45,0x05,0x43,0x00,0x27,0x03,0x28,0x00,0x33,0x04,0x49,0x00,0x45,0x03,0x94,0x00,0x12,0x04,0xa7,0x00,0x35,0x04,0x22,0x00,0x11,0x06,0x6d,0x00,0x08,0x04,0x22,0x00,0x1c,0x04,0x9e,0x00,0x32,0x03,0xca,0x00,0x32,0x03,0xf6,0x00,0x87,0x02,0x3b,0x00,0x9c,0x04,0x2d,0x00,0x33,0x05,0xc5,0x00,0x07,0x04,0x00,0x01,0x00,0x03,0x2f,0x00,0x16,0x03,0xf6,0x00,0x57,0x03,0x14,0x00,0x34,0x02,0xa2,0x00,0x3c,0x04,0x73,0x00,0x28,0x04,0x73,0x00,0x20,0x04,0x00,0x00,0xd3,0x02,0xc4,0x00,0x9e,0x04,0x00,0x01,0x58,0x04,0x73,0x00,0xbd,0x06,0xac,0x00,0x1b,0x06,0x52,0x00,0x1a,0x06,0xac,0x00,0x20,0x00,0x00,0x00,0x03,0x00,0x00,0x00,0x03,0x00,0x00,0x00,0x1c,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0xa0,0x00,0x03,0x00,0x01,0x00,0x00,0x00,0x1c,0x00,0x04,0x00,0x84,0x00,0x00,0x00,0x1a,0x00,0x10,0x00,0x03,0x00,0x0a,0x00,0x7a,0x00,0x7e,0x00,0xa3,0x00,0xa8,0x00,0xaa,0x00,0xad,0x00,0xb0,0x00,0xb4,0x00,0xb9,0x00,0xbe,0x03,0x7e,0x22,0x19,0xff,0xff,0x00,0x00,0x00,0x20,0x00,0x7e,0x00,0xa0,0x00,0xa8,0x00,0xaa,0x00,0xac,0x00,0xaf,0x00,0xb2,0x00,0xb7,0x00,0xbc,0x03,0x7e,0x22,0x19,0xff,0xff,0xff,0xe3,0xff,0xe0,0x00,0x00,0xff,0xba,0xff,0xb9,0x00,0x00,0xff,0xb6,0xff,0xb5,0xff,0xb3,0xff,0xb1,0xfc,0xa0,0xde,0x51,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x16,0x00,0x00,0x00,0x00,0x00,0x18,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x03,0x00,0x5f,0x00,0x60,0x00,0x61,0x00,0x64,0x00,0x10,0x00,0x06,0x02,0x04,0x00,0x00,0x00,0x00,0x00,0xfd,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x01,0x00,0x02,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x02,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x03,0x00,0x04,0x00,0x05,0x00,0x06,0x00,0x07,0x00,0x08,0x00,0x09,0x00,0x0a,0x00,0x0b,0x00,0x0c,0x00,0x0d,0x00,0x0e,0x00,0x0f,0x00,0x10,0x00,0x11,0x00,0x12,0x00,0x13,0x00,0x14,0x00,0x15,0x00,0x16,0x00,0x17,0x00,0x18,0x00,0x19,0x00,0x1a,0x00,0x1b,0x00,0x1c,0x00,0x1d,0x00,0x1e,0x00,0x1f,0x00,0x20,0x00,0x21,0x00,0x22,0x00,0x23,0x00,0x24,0x00,0x25,0x00,0x26,0x00,0x27,0x00,0x28,0x00,0x29,0x00,0x2a,0x00,0x2b,0x00,0x2c,0x00,0x2d,0x00,0x2e,0x00,0x2f,0x00,0x30,0x00,0x31,0x00,0x32,0x00,0x33,0x00,0x34,0x00,0x35,0x00,0x36,0x00,0x37,0x00,0x38,0x00,0x39,0x00,0x3a,0x00,0x3b,0x00,0x3c,0x00,0x3d,0x00,0x3e,0x00,0x3f,0x00,0x40,0x00,0x41,0x00,0x42,0x00,0x43,0x00,0x44,0x00,0x45,0x00,0x46,0x00,0x47,0x00,0x48,0x00,0x49,0x00,0x4a,0x00,0x4b,0x00,0x4c,0x00,0x4d,0x00,0x4e,0x00,0x4f,0x00,0x50,0x00,0x51,0x00,0x52,0x00,0x53,0x00,0x54,0x00,0x55,0x00,0x56,0x00,0x57,0x00,0x58,0x00,0x59,0x00,0x5a,0x00,0x5b,0x00,0x5c,0x00,0x5d,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x5e,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x66,0x00,0x60,0x00,0x61,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x69,0x00,0x62,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x63,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x5f,0x00,0x64,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x03,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x6a,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x65,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x6b,0x00,0x00,0x00,0x56,0x00,0x56,0x00,0x56,0x00,0x56,0x00,0x7c,0x00,0xa4,0x01,0x34,0x01,0xda,0x02,0x4a,0x02,0xa6,0x02,0xbe,0x02,0xea,0x03,0x16,0x03,0x58,0x03,0x80,0x03,0x98,0x03,0xb0,0x03,0xc2,0x03,0xe0,0x04,0x12,0x04,0x38,0x04,0x76,0x04,0xc0,0x04,0xfa,0x05,0x48,0x05,0x8c,0x05,0xbc,0x06,0x0a,0x06,0x48,0x06,0x68,0x06,0x8c,0x06,0xb4,0x06,0xdc,0x07,0x04,0x07,0x40,0x07,0xb2,0x07,0xea,0x08,0x3c,0x08,0x72,0x08,0xae,0x08,0xde,0x09,0x08,0x09,0x52,0x09,0x8e,0x09,0xb0,0x09,0xea,0x0a,0x2c,0x0a,0x52,0x0a,0x8a,0x0a,0xb6,0x0b,0x04,0x0b,0x3c,0x0b,0x98,0x0b,0xda,0x0c,0x1c,0x0c,0x3a,0x0c,0x6e,0x0c,0x96,0x0c,0xe0,0x0d,0x1c,0x0d,0x48,0x0d,0x76,0x0d,0x98,0x0d,0xb6,0x0d,0xd8,0x0d,0xd8,0x0d,0xee,0x0e,0x0c,0x0e,0x54,0x0e,0x8e,0x0e,0xc0,0x0f,0x00,0x0f,0x3c,0x0f,0x70,0x0f,0xbc,0x0f,0xf0,0x10,0x1e,0x10,0x52,0x10,0x88,0x10,0xaa,0x10,0xfa,0x11,0x30,0x11,0x6a,0x11,0xa8,0x11,0xee,0x12,0x1a,0x12,0x56,0x12,0x90,0x12,0xc6,0x12,0xf2,0x13,0x3a,0x13,0x78,0x13,0xba,0x13,0xe4,0x14,0x0e,0x14,0x18,0x14,0x74,0x14,0xd0,0x14,0xee,0x15,0x00,0x15,0x12,0x15,0x30,0x15,0x56,0x15,0x94,0x15,0xde,0x15,0xfa,0x16,0x0e,0x16,0x36,0x16,0x5c,0x16,0xc4,0x17,0x2e,0x17,0xb6,0x00,0x00,0x00,0x04,0x00,0x64,0x00,0x00,0x03,0x9c,0x05,0x9a,0x00,0x03,0x00,0x07,0x00,0x24,0x00,0x38,0x00,0x00,0x33,0x11,0x21,0x11,0x25,0x21,0x11,0x21,0x17,0x36,0x37,0x36,0x33,0x32,0x16,0x15,0x14,0x06,0x07,0x0e,0x01,0x15,0x14,0x17,0x23,0x26,0x35,0x34,0x12,0x35,0x34,0x26,0x23,0x22,0x07,0x06,0x07,0x13,0x37,0x36,0x33,0x32,0x1f,0x01,0x16,0x15,0x14,0x0f,0x01,0x06,0x23,0x22,0x2f,0x01,0x26,0x35,0x34,0x64,0x03,0x38,0xfc,0xfa,0x02,0xd4,0xfd,0x2c,0xaf,0x1f,0x1b,0x35,0x3b,0x5c,0x70,0x2e,0x40,0x3f,0x48,0x18,0x20,0x23,0xa3,0x42,0x3a,0x26,0x1f,0x1a,0x1e,0x40,0x39,0x0b,0x09,0x0a,0x0c,0x38,0x09,0x0a,0x38,0x0e,0x07,0x0b,0x09,0x3d,0x07,0x05,0x9a,0xfa,0x66,0x32,0x05,0x36,0xec,0x1c,0x0f,0x1e,0x5f,0x50,0x31,0x63,0x50,0x50,0x68,0x2f,0x26,0x5f,0x61,0x33,0x4c,0x01,0x1c,0x4b,0x39,0x42,0x11,0x0f,0x19,0xfc,0xff,0x3a,0x0a,0x0b,0x3c,0x0b,0x09,0x0b,0x0b,0x3e,0x0e,0x0a,0x47,0x09,0x09,0x0a,0x00,0x02,0x00,0xce,0xff,0xfe,0x01,0xd2,0x06,0xc1,0x00,0x0b,0x00,0x13,0x00,0x00,0x01,0x26,0x35,0x02,0x27,0x36,0x33,0x16,0x17,0x14,0x03,0x14,0x02,0x37,0x32,0x17,0x14,0x07,0x26,0x27,0x01,0x3e,0x65,0x07,0x01,0x01,0x70,0x70,0x05,0x0a,0xde,0x76,0x83,0x0a,0x7b,0x7f,0x0a,0x02,0x03,0x19,0x5c,0x03,0x82,0x4c,0x7b,0x02,0x7c,0x50,0xfc,0x7e,0x5d,0xfe,0xeb,0x0a,0x7f,0x89,0x03,0x01,0x7a,0x00,0x00,0x02,0x00,0x64,0x05,0x0b,0x02,0x58,0x07,0x41,0x00,0x09,0x00,0x13,0x00,0x00,0x00,0x17,0x03,0x06,0x07,0x26,0x35,0x03,0x36,0x33,0x04,0x17,0x03,0x06,0x07,0x26,0x35,0x03,0x36,0x33,0x01,0x23,0x09,0x0d,0x01,0x57,0x57,0x0c,0x14,0x52,0x01,0x85,0x09,0x0d,0x01,0x57,0x57,0x0c,0x14,0x52,0x07,0x3d,0x51,0xfe,0x8a,0x6a,0x01,0x01,0x6f,0x01,0x75,0x51,0x04,0x51,0xfe,0x8a,0x6a,0x01,0x01,0x6f,0x01,0x75,0x51,0x00,0x00,0x02,0x00,0x41,0xff,0xf8,0x04,0xbb,0x06,0x5c,0x00,0x09,0x00,0x5a,0x00,0x00,0x01,0x06,0x07,0x06,0x07,0x36,0x37,0x13,0x36,0x37,0x05,0x07,0x26,0x27,0x36,0x37,0x32,0x37,0x32,0x37,0x36,0x37,0x36,0x33,0x16,0x17,0x06,0x07,0x36,0x37,0x36,0x37,0x36,0x33,0x16,0x17,0x06,0x07,0x16,0x33,0x16,0x17,0x06,0x07,0x06,0x07,0x26,0x27,0x26,0x27,0x06,0x07,0x06,0x07,0x16,0x33,0x16,0x17,0x06,0x07,0x06,0x07,0x26,0x27,0x26,0x23,0x02,0x07,0x26,0x35,0x36,0x13,0x07,0x02,0x07,0x26,0x35,0x34,0x13,0x07,0x26,0x27,0x36,0x37,0x32,0x37,0x36,0x37,0x13,0x36,0x37,0x02,0x5b,0x16,0x1b,0x17,0x16,0x4b,0x5b,0x5c,0x06,0x06,0xfe,0x5d,0x6a,0x46,0x04,0x0e,0x3d,0x23,0x68,0x1f,0x26,0x25,0x16,0x22,0x36,0x45,0x08,0x02,0x2f,0x50,0x61,0x23,0x16,0x22,0x35,0x45,0x08,0x02,0x2e,0x77,0x1d,0x3d,0x0e,0x02,0x1c,0x0c,0x1d,0x0f,0x10,0x73,0x28,0x16,0x1d,0x16,0x15,0x7a,0x22,0x3d,0x0e,0x02,0x11,0x08,0x27,0x13,0x14,0x76,0x2e,0x75,0x5f,0x52,0x01,0x5f,0x9a,0x74,0x5e,0x51,0x5b,0x83,0x46,0x04,0x0e,0x3d,0x29,0x8d,0x01,0x01,0x5e,0x05,0x05,0x04,0x37,0x68,0x7e,0x75,0x65,0x01,0x02,0x01,0x89,0x1b,0x1b,0x0c,0x08,0x0c,0x51,0x50,0x04,0x02,0x01,0xb2,0x98,0x39,0x04,0x60,0x33,0xe8,0x02,0x02,0xaa,0x93,0x39,0x03,0x61,0x32,0xe2,0x04,0x04,0x50,0x32,0x18,0x12,0x06,0x04,0x03,0x0f,0x01,0x6b,0x85,0x70,0x62,0x03,0x04,0x50,0x26,0x17,0x1f,0x07,0x05,0x03,0x0e,0xfe,0x23,0x01,0x03,0x4c,0x4b,0x01,0x41,0x03,0xfe,0x2e,0x01,0x02,0x4c,0x4b,0x01,0x33,0x09,0x0b,0x52,0x4f,0x04,0x03,0x03,0x04,0x01,0x8d,0x16,0x15,0x00,0x00,0x05,0x00,0x45,0xfe,0xc4,0x04,0xa5,0x07,0x56,0x00,0x44,0x00,0x4b,0x00,0x52,0x00,0x5c,0x00,0x67,0x00,0x00,0x01,0x36,0x37,0x32,0x17,0x11,0x36,0x37,0x16,0x17,0x11,0x16,0x17,0x16,0x15,0x14,0x07,0x06,0x23,0x22,0x27,0x26,0x27,0x11,0x16,0x17,0x16,0x15,0x02,0x05,0x11,0x06,0x07,0x26,0x27,0x11,0x06,0x07,0x23,0x26,0x27,0x11,0x06,0x07,0x26,0x27,0x11,0x26,0x27,0x26,0x35,0x37,0x36,0x33,0x32,0x17,0x16,0x17,0x11,0x24,0x03,0x37,0x12,0x25,0x11,0x36,0x37,0x16,0x17,0x01,0x36,0x37,0x36,0x35,0x34,0x27,0x01,0x06,0x07,0x06,0x15,0x14,0x17,0x05,0x26,0x27,0x26,0x27,0x11,0x16,0x17,0x36,0x37,0x11,0x26,0x2b,0x01,0x06,0x07,0x11,0x16,0x17,0x16,0x17,0x02,0x2a,0x1c,0x1e,0x45,0x31,0x01,0x47,0x47,0x01,0x66,0x3c,0x62,0x08,0x11,0x1d,0x2e,0x4a,0x22,0x34,0x91,0x3c,0x6e,0x0b,0xfe,0xd0,0x01,0x47,0x47,0x01,0x14,0x21,0x49,0x19,0x19,0x01,0x3d,0x51,0x01,0x55,0x5c,0xa4,0x11,0x14,0x15,0x44,0x51,0x39,0x4d,0xfe,0xe5,0x14,0x02,0x18,0x01,0x15,0x01,0x51,0x3d,0x01,0x01,0x40,0x90,0x0e,0x01,0x9f,0xfe,0x30,0x83,0x03,0x05,0x8b,0x01,0x40,0x3d,0x5a,0x0d,0x0c,0x26,0x2a,0x39,0x27,0x2e,0x40,0x03,0x21,0x1e,0x12,0x14,0x50,0x3a,0x06,0x0f,0x02,0x02,0x09,0x01,0x09,0x42,0x01,0x01,0x43,0xfe,0xd9,0x22,0x3f,0x69,0x48,0x14,0x12,0x20,0x54,0x27,0x1c,0xfe,0x69,0x27,0x49,0x86,0xd4,0xfe,0xcc,0x5d,0xfe,0xcd,0x40,0x01,0x01,0x44,0x01,0x13,0x04,0x03,0x01,0x03,0xfe,0xec,0x40,0x01,0x01,0x44,0x01,0x2f,0x29,0x5a,0x9f,0xae,0x17,0x0e,0x96,0x68,0x35,0x02,0x15,0x41,0x01,0x14,0x2b,0x01,0x1e,0x4c,0x01,0x1a,0x42,0x01,0x01,0x43,0xf9,0xe3,0x3f,0x8a,0x09,0x09,0xa3,0x4b,0x02,0x83,0x3c,0x7a,0x14,0x12,0x6c,0x28,0xe9,0x10,0x04,0x01,0x01,0xfd,0xcf,0x07,0x03,0x03,0x09,0x04,0x90,0x0e,0x04,0x06,0xfe,0x5b,0x02,0x01,0x04,0x0a,0x00,0x00,0x05,0x00,0x20,0xff,0xeb,0x06,0x76,0x06,0x25,0x00,0x0d,0x00,0x19,0x00,0x27,0x00,0x33,0x00,0x41,0x00,0x00,0x01,0x17,0x1e,0x01,0x17,0x14,0x06,0x07,0x27,0x2e,0x01,0x27,0x3e,0x01,0x03,0x16,0x1f,0x01,0x36,0x3f,0x01,0x34,0x26,0x27,0x23,0x06,0x01,0x17,0x1e,0x01,0x17,0x14,0x06,0x07,0x27,0x2e,0x01,0x27,0x3e,0x01,0x03,0x16,0x1f,0x01,0x36,0x3f,0x01,0x34,0x26,0x27,0x23,0x06,0x00,0x37,0x32,0x17,0x14,0x07,0x01,0x06,0x07,0x26,0x27,0x36,0x37,0x01,0x01,0x82,0x2e,0x7d,0xe1,0x1a,0xc0,0xb8,0x22,0xa1,0xc8,0x05,0x09,0xae,0x28,0x0c,0xc4,0x2b,0xb3,0x2a,0x05,0x93,0x63,0x1c,0xb4,0x04,0x0a,0x2d,0x7e,0xe1,0x1a,0xc1,0xb8,0x21,0xa1,0xc8,0x05,0x08,0xae,0x28,0x0d,0xc4,0x2a,0xb4,0x2a,0x05,0x93,0x63,0x1c,0xb4,0x01,0x96,0x3d,0x27,0x13,0x32,0xfb,0x52,0x44,0x39,0x32,0x0b,0x07,0x3e,0x04,0xbd,0x06,0x25,0x02,0x08,0xbc,0xbd,0xb6,0xc9,0x0d,0x05,0x11,0xd3,0xc1,0x95,0xc6,0xfe,0x99,0xd3,0x3a,0x06,0x12,0xac,0x1b,0x77,0x99,0x0a,0x18,0xfd,0xa7,0x01,0x08,0xbd,0xbd,0xb6,0xc9,0x0c,0x04,0x11,0xd3,0xc1,0x95,0xc7,0xfe,0x98,0xd3,0x39,0x07,0x12,0xac,0x1c,0x77,0x99,0x09,0x17,0x03,0x94,0x03,0x3d,0x43,0x2a,0xfa,0xd1,0x45,0x09,0x09,0x50,0x3d,0x34,0x05,0x37,0x00,0x03,0x00,0x92,0xff,0xf7,0x06,0xa0,0x07,0x4a,0x00,0x21,0x00,0x29,0x00,0x31,0x00,0x00,0x24,0x17,0x06,0x07,0x26,0x2f,0x01,0x06,0x05,0x23,0x24,0x03,0x35,0x12,0x01,0x26,0x35,0x36,0x25,0x33,0x04,0x13,0x06,0x07,0x16,0x13,0x36,0x13,0x34,0x37,0x16,0x15,0x02,0x07,0x01,0x06,0x07,0x16,0x17,0x36,0x37,0x34,0x03,0x04,0x03,0x12,0x05,0x36,0x37,0x02,0x06,0x46,0x14,0x03,0x70,0x50,0x2b,0x2a,0xc3,0xfe,0xcf,0x5b,0xfd,0xb4,0x15,0x11,0x01,0x89,0xd0,0x1f,0x01,0x51,0x4c,0x01,0x32,0x09,0x0a,0xbc,0xfe,0xec,0x44,0x22,0x63,0x60,0x15,0x9e,0xfc,0xf6,0xaa,0x05,0x2f,0x85,0x69,0x3b,0xae,0xfe,0x9b,0x0f,0x16,0x01,0x95,0xef,0xde,0xb2,0xb5,0x4f,0x6d,0x01,0x15,0x5f,0x61,0xbc,0x1a,0x12,0x01,0xee,0x52,0x01,0x67,0x01,0x23,0x82,0xf1,0xf6,0x0e,0x0c,0xfe,0xd3,0xc5,0x9b,0xaf,0xfe,0x4d,0x6f,0x01,0x18,0x76,0x04,0x04,0x86,0xfe,0xa0,0xfe,0x05,0x1b,0x03,0x83,0x82,0x32,0x28,0x88,0x8a,0xfd,0xaa,0xdc,0xfe,0xca,0xfe,0xb9,0x05,0x01,0xbf,0x01,0x9a,0x00,0x00,0x00,0x01,0x00,0x64,0x05,0x0b,0x01,0x2c,0x07,0x41,0x00,0x09,0x00,0x00,0x00,0x17,0x03,0x06,0x07,0x26,0x35,0x03,0x36,0x33,0x01,0x23,0x09,0x0d,0x01,0x57,0x57,0x0c,0x14,0x52,0x07,0x3d,0x51,0xfe,0x8a,0x6a,0x01,0x01,0x6f,0x01,0x75,0x51,0x00,0x00,0x00,0x01,0x00,0x7d,0xfe,0x74,0x02,0x89,0x08,0x05,0x00,0x15,0x00,0x00,0x00,0x37,0x16,0x17,0x06,0x07,0x02,0x03,0x10,0x13,0x16,0x17,0x06,0x07,0x22,0x27,0x26,0x27,0x02,0x03,0x12,0x13,0x01,0xa6,0x7c,0x53,0x09,0x12,0x5c,0xc0,0x0d,0xc4,0x5b,0x27,0x01,0x4f,0x5a,0x30,0x3e,0x32,0xc1,0x01,0x0c,0xcb,0x08,0x01,0x04,0x15,0x65,0x62,0x8f,0xfe,0xd9,0xfe,0x17,0xfe,0x1d,0xfe,0x6a,0xa6,0x7c,0x73,0x08,0x3e,0x55,0x83,0x02,0x0a,0x01,0xdb,0x02,0x06,0x01,0xa3,0x00,0x01,0x00,0x51,0xfe,0x74,0x02,0x62,0x08,0x0a,0x00,0x15,0x00,0x00,0x12,0x27,0x34,0x37,0x16,0x17,0x12,0x13,0x02,0x03,0x06,0x07,0x06,0x07,0x22,0x27,0x36,0x37,0x12,0x13,0x02,0x03,0x81,0x1a,0x62,0x5b,0x4d,0xf0,0x01,0x01,0xb4,0x46,0x44,0x2e,0x44,0x59,0x07,0x0a,0x66,0xda,0x02,0x0a,0xb5,0x07,0x0e,0x7f,0x73,0x0a,0x0a,0xab,0xfe,0x5f,0xfd,0xa6,0xfe,0x1e,0xfe,0x35,0xaf,0x4d,0x35,0x08,0x6b,0x55,0x8a,0x01,0xbf,0x01,0xf8,0x01,0xce,0x01,0x50,0x00,0x00,0x01,0x00,0x4c,0x03,0xe6,0x02,0xe1,0x06,0xf3,0x00,0x27,0x00,0x00,0x01,0x26,0x35,0x36,0x33,0x32,0x17,0x14,0x07,0x36,0x37,0x16,0x15,0x06,0x07,0x16,0x17,0x06,0x07,0x26,0x27,0x16,0x15,0x06,0x07,0x26,0x27,0x36,0x37,0x06,0x07,0x26,0x27,0x36,0x37,0x26,0x27,0x36,0x37,0x16,0x01,0x64,0x1b,0x1c,0x30,0x30,0x1d,0x18,0x74,0x74,0x2c,0x21,0xab,0xc8,0x07,0x07,0x2c,0x50,0x88,0x12,0x09,0x40,0x49,0x09,0x01,0x12,0x7b,0x43,0x45,0x04,0x05,0xc7,0xbf,0x1a,0x01,0x3a,0x57,0x05,0xd9,0x84,0x4f,0x47,0x48,0x47,0x90,0xae,0x02,0x0d,0x3f,0x6c,0x50,0x53,0x5c,0x33,0x0e,0x08,0x76,0x7e,0x5b,0x48,0x03,0x0f,0x55,0x41,0x83,0x75,0x07,0x06,0x3d,0x43,0x69,0x4a,0x6e,0x3e,0x10,0x01,0x00,0x00,0x00,0x01,0x00,0xc0,0x00,0xc7,0x03,0xf3,0x03,0xed,0x00,0x17,0x00,0x00,0x01,0x33,0x16,0x17,0x06,0x07,0x23,0x15,0x06,0x07,0x26,0x3d,0x01,0x23,0x26,0x27,0x36,0x3b,0x01,0x35,0x36,0x37,0x16,0x17,0x02,0xc7,0x9b,0x84,0x0d,0x07,0x82,0xa2,0x06,0x68,0x5c,0xaf,0x8b,0x04,0x08,0x89,0xac,0x01,0x5d,0x60,0x0c,0x02,0xc9,0x01,0x5d,0x60,0x0c,0xab,0x89,0x04,0x08,0x86,0xa9,0x06,0x68,0x5c,0x97,0x81,0x0d,0x07,0x80,0x00,0x00,0x01,0x00,0x9e,0xfe,0xf1,0x01,0x66,0x00,0xe1,0x00,0x09,0x00,0x00,0x24,0x17,0x03,0x06,0x07,0x26,0x35,0x03,0x36,0x33,0x01,0x5d,0x09,0x0d,0x01,0x57,0x57,0x0c,0x14,0x52,0xdd,0x51,0xfe,0xd0,0x6a,0x01,0x01,0x6f,0x01,0x2f,0x51,0x00,0x00,0x00,0x00,0x01,0x00,0x14,0x02,0x63,0x02,0xe4,0x03,0x2e,0x00,0x09,0x00,0x00,0x00,0x17,0x06,0x07,0x05,0x26,0x27,0x36,0x33,0x25,0x02,0xd8,0x0c,0x06,0x72,0xfe,0x26,0x7a,0x04,0x07,0x78,0x01,0xd2,0x03,0x2d,0x5d,0x60,0x0c,0x01,0x06,0x68,0x5c,0x01,0x00,0x00,0x01,0x00,0x9e,0xff,0xfe,0x01,0xa2,0x01,0x09,0x00,0x07,0x00,0x00,0x36,0x37,0x32,0x17,0x14,0x07,0x26,0x27,0x9f,0x76,0x83,0x0a,0x7b,0x7f,0x0a,0xff,0x0a,0x7f,0x89,0x03,0x01,0x7a,0x00,0x01,0xff,0xf7,0xff,0xe0,0x03,0x38,0x07,0x4f,0x00,0x0d,0x00,0x00,0x01,0x16,0x17,0x06,0x07,0x01,0x06,0x23,0x26,0x27,0x34,0x37,0x01,0x36,0x02,0xf5,0x42,0x01,0x06,0x1c,0xfd,0x80,0x1f,0x3a,0x40,0x06,0x25,0x02,0x80,0x13,0x07,0x4f,0x05,0x61,0x3c,0x36,0xf9,0xbe,0x55,0x04,0x44,0x2c,0x56,0x06,0x43,0x58,0x00,0x02,0x00,0x0d,0xff,0xf1,0x04,0x64,0x05,0xca,0x00,0x0b,0x00,0x15,0x00,0x00,0x01,0x17,0x04,0x13,0x17,0x02,0x05,0x27,0x24,0x03,0x27,0x12,0x13,0x12,0x05,0x20,0x13,0x27,0x02,0x25,0x04,0x03,0x02,0x38,0x44,0x01,0x92,0x50,0x06,0x22,0xfd,0xdb,0x43,0xfe,0x77,0x36,0x0e,0x0f,0xad,0x11,0x01,0x11,0x01,0x9e,0x24,0x05,0x34,0xfe,0xd7,0xfe,0xb4,0x3a,0x05,0xca,0x03,0x37,0xfd,0xf2,0x88,0xfd,0x0e,0x17,0x03,0x64,0x01,0xae,0x85,0x03,0x18,0xfc,0xee,0xfe,0x67,0x4a,0x02,0x33,0x6b,0x01,0xb4,0x12,0x15,0xfd,0xe6,0x00,0x00,0x01,0x00,0xa9,0x00,0x00,0x03,0x13,0x05,0xc1,0x00,0x12,0x00,0x00,0x00,0x17,0x02,0x03,0x06,0x23,0x26,0x27,0x12,0x11,0x06,0x07,0x26,0x27,0x34,0x3f,0x01,0x36,0x33,0x02,0xfe,0x15,0x05,0x15,0x09,0x5e,0x57,0x11,0x23,0xe3,0x66,0x48,0x13,0x2f,0xe4,0x8b,0x59,0x05,0xb7,0x40,0xfe,0x08,0xfc,0xc4,0x43,0x03,0x3e,0x03,0x3d,0x01,0x51,0xf9,0x0c,0x07,0x3d,0x48,0x25,0xba,0x8c,0x00,0x00,0x00,0x00,0x01,0x00,0x28,0xff,0xf6,0x04,0x48,0x05,0xb7,0x00,0x20,0x00,0x00,0x01,0x04,0x13,0x14,0x02,0x05,0x25,0x32,0x16,0x17,0x14,0x23,0x26,0x27,0x04,0x07,0x26,0x35,0x36,0x25,0x24,0x11,0x02,0x25,0x04,0x03,0x06,0x23,0x22,0x27,0x37,0x12,0x25,0x02,0x5c,0x01,0x9b,0x35,0xfa,0xfe,0x7c,0x01,0x0e,0x91,0xf5,0x06,0x6f,0x44,0xd5,0xfe,0x69,0x6f,0x67,0x01,0x01,0x83,0x01,0x92,0x18,0xfe,0xed,0xfe,0xea,0x3a,0x0a,0x5d,0x5e,0x01,0x02,0x44,0x01,0x9a,0x05,0xb7,0x2b,0xfe,0x62,0xe5,0xfe,0xb2,0xe9,0x12,0x30,0x62,0x57,0x19,0x0c,0x11,0x19,0x0a,0x61,0x7e,0xfc,0xe7,0x01,0x1f,0x01,0x09,0x19,0x0a,0xfe,0xf8,0x74,0x6a,0x1f,0x01,0x83,0x2e,0x00,0x00,0x00,0x01,0x00,0x20,0xff,0xf7,0x04,0x57,0x05,0xc5,0x00,0x27,0x00,0x00,0x01,0x04,0x1f,0x01,0x06,0x07,0x04,0x13,0x02,0x05,0x24,0x03,0x36,0x33,0x32,0x12,0x17,0x24,0x37,0x02,0x25,0x06,0x07,0x26,0x35,0x36,0x37,0x36,0x35,0x26,0x27,0x04,0x07,0x14,0x07,0x26,0x27,0x37,0x12,0x25,0x02,0x69,0x01,0x1c,0x3d,0x0a,0x08,0x87,0x01,0x15,0x05,0x33,0xfe,0x16,0xfe,0x00,0x1a,0x0e,0x54,0x42,0x62,0xfb,0x01,0x49,0x23,0x13,0xfe,0xfd,0x5e,0x6c,0x61,0x0b,0xd0,0xcb,0x11,0x86,0xfe,0xbd,0x32,0x5e,0x4c,0x09,0x01,0x49,0x01,0x8f,0x05,0xc5,0x18,0xee,0x3c,0x9e,0x74,0x55,0xfe,0xab,0xfe,0x5d,0x2d,0x04,0x01,0x98,0x47,0xfe,0xfe,0x14,0x0e,0xfb,0x01,0x14,0x0e,0x07,0x07,0x14,0x54,0x5d,0x19,0x18,0xc1,0x72,0x07,0x07,0xc7,0x46,0x0a,0x14,0x55,0x32,0x01,0x20,0x15,0x00,0x00,0x00,0x00,0x02,0x00,0x00,0xff,0xf6,0x04,0x6a,0x05,0xc8,0x00,0x17,0x00,0x1d,0x00,0x00,0x01,0x32,0x17,0x02,0x03,0x37,0x16,0x17,0x06,0x23,0x27,0x13,0x06,0x23,0x26,0x27,0x37,0x04,0x05,0x26,0x3d,0x01,0x12,0x00,0x17,0x00,0x03,0x36,0x37,0x12,0x02,0xe4,0x80,0x14,0x03,0x23,0xa4,0x60,0x14,0x0b,0x49,0xc4,0x05,0x10,0x56,0x54,0x0a,0x09,0xfe,0xe4,0xfe,0xe3,0x63,0x25,0x02,0x74,0x2b,0xfe,0x18,0x09,0xd4,0xf8,0x22,0x05,0xc8,0x6b,0xfe,0x7b,0xfe,0x1f,0x0b,0x09,0x5e,0x6c,0x08,0xff,0x00,0x41,0x07,0x5d,0xd4,0x02,0x35,0x0f,0x88,0x2a,0x01,0x2d,0x02,0xe3,0xed,0xfe,0x00,0xfe,0xe9,0x2d,0x02,0x01,0xf1,0x00,0x00,0x01,0x00,0x35,0xff,0xf2,0x04,0x46,0x05,0xc1,0x00,0x2c,0x00,0x00,0x01,0x36,0x37,0x32,0x17,0x0e,0x01,0x07,0x25,0x06,0x07,0x17,0x3e,0x01,0x37,0x16,0x12,0x1d,0x01,0x02,0x05,0x07,0x22,0x00,0x35,0x36,0x37,0x32,0x17,0x16,0x17,0x36,0x13,0x37,0x02,0x27,0x0e,0x01,0x07,0x22,0x27,0x12,0x3f,0x01,0x16,0x02,0x52,0x8f,0x7a,0x58,0x08,0x01,0x8b,0xd5,0xfe,0xf9,0x56,0x02,0x0d,0x52,0xc7,0x87,0xe0,0xbe,0x28,0xfe,0x97,0x87,0xd2,0xfe,0xd9,0x07,0x4a,0x49,0x35,0x6b,0xe9,0xff,0x2f,0x04,0x0f,0xe9,0x71,0xe8,0x5c,0x8a,0x14,0x22,0x93,0x21,0x6d,0x05,0xa5,0x08,0x14,0x52,0x51,0x2c,0x06,0x05,0x8d,0x6f,0x0f,0x0c,0x37,0x0a,0x06,0xfe,0xdc,0xba,0x4d,0xfe,0x23,0x2d,0x06,0x01,0x03,0x76,0x41,0x0a,0x59,0xa6,0x01,0x0a,0x01,0x2c,0x69,0x01,0x0c,0x0f,0x0d,0x3f,0x04,0xae,0x01,0x3a,0xaa,0x07,0x10,0x00,0x00,0x00,0x00,0x02,0x00,0x0a,0x00,0x00,0x04,0x66,0x05,0xb8,0x00,0x19,0x00,0x23,0x00,0x00,0x01,0x17,0x16,0x17,0x06,0x07,0x2e,0x01,0x27,0x06,0x02,0x07,0x36,0x37,0x33,0x04,0x13,0x07,0x02,0x05,0x24,0x03,0x35,0x10,0x37,0x36,0x03,0x15,0x12,0x05,0x33,0x24,0x13,0x10,0x25,0x04,0x02,0x40,0x3c,0xf7,0x11,0x0c,0x55,0x5a,0x41,0x41,0x94,0xdc,0x0e,0x8b,0xf2,0x21,0x01,0xd5,0x2a,0x01,0x1f,0xfe,0x1e,0xfd,0xb8,0x12,0x96,0xcb,0x9d,0x22,0x01,0x53,0x26,0x01,0x36,0x0a,0xfe,0xc3,0xfe,0xbb,0x05,0xb8,0x01,0x20,0x74,0x52,0x06,0x0a,0x24,0x10,0x0e,0xfe,0xdf,0x9a,0xa8,0x12,0x1f,0xfe,0x70,0x6b,0xfe,0x76,0x56,0x06,0x02,0x55,0x4a,0x01,0x39,0xdd,0xfc,0xfc,0x6c,0x37,0xfe,0xdd,0x0a,0x4c,0x01,0x0f,0x01,0x05,0x26,0x25,0x00,0x01,0x00,0x1a,0xff,0xfb,0x04,0x4d,0x05,0xc0,0x00,0x19,0x00,0x00,0x01,0x16,0x17,0x14,0x07,0x00,0x03,0x15,0x06,0x23,0x22,0x35,0x37,0x12,0x25,0x06,0x07,0x27,0x26,0x27,0x34,0x37,0x16,0x17,0x36,0x24,0x03,0xc4,0x7f,0x0a,0x3b,0xfe,0x42,0x10,0x12,0x5a,0x69,0x01,0x4e,0x01,0x3a,0x77,0xe7,0x91,0xe7,0x08,0x66,0xcc,0x70,0x5e,0x01,0x39,0x05,0xc0,0x0a,0x53,0x3f,0x28,0xfe,0xc5,0xfd,0xa6,0xf0,0x7c,0x85,0xf0,0x02,0x91,0xfc,0x2b,0x0d,0x0d,0x14,0x63,0x5c,0x0d,0x21,0x04,0x06,0x2d,0x00,0x00,0x00,0x03,0x00,0x11,0xff,0xef,0x04,0x61,0x05,0xd6,0x00,0x15,0x00,0x1d,0x00,0x27,0x00,0x00,0x01,0x33,0x04,0x13,0x17,0x06,0x07,0x04,0x13,0x15,0x02,0x05,0x27,0x24,0x03,0x35,0x12,0x37,0x26,0x27,0x37,0x12,0x13,0x16,0x17,0x36,0x37,0x26,0x27,0x06,0x02,0x07,0x16,0x05,0x37,0x24,0x13,0x26,0x25,0x07,0x02,0x2d,0x2a,0x01,0x23,0x3b,0x01,0x09,0x7b,0x01,0x16,0x19,0x25,0xfe,0x13,0x60,0xfe,0x4d,0x2b,0x10,0xcd,0x67,0x0a,0x04,0x2d,0x92,0x05,0xbd,0xe7,0x11,0x1a,0x8c,0xfb,0x87,0x07,0x01,0x01,0x46,0x34,0x01,0x51,0x06,0x1b,0xfe,0x9d,0x51,0x05,0xd6,0x01,0xfe,0xff,0x2d,0xd0,0x55,0x3e,0xfe,0xeb,0x37,0xfe,0x11,0x1a,0x02,0x16,0x01,0x6d,0x3c,0x01,0x17,0x8a,0x66,0x98,0x29,0x01,0x33,0xfe,0xb8,0xae,0x04,0x29,0xc1,0x8c,0x08,0x0c,0xfd,0x6a,0xf5,0xc9,0x2a,0x01,0x32,0x01,0x34,0xd4,0x11,0x0d,0x00,0x00,0x00,0x00,0x02,0x00,0x21,0xff,0xfe,0x04,0x53,0x05,0xc1,0x00,0x13,0x00,0x1e,0x00,0x00,0x01,0x04,0x13,0x02,0x05,0x27,0x26,0x35,0x34,0x24,0x00,0x13,0x27,0x02,0x05,0x24,0x03,0x10,0x37,0x36,0x03,0x16,0x17,0x20,0x13,0x27,0x2e,0x01,0x23,0x07,0x06,0x02,0x08,0x02,0x26,0x25,0x20,0xfd,0x3b,0x4d,0x42,0x01,0xa3,0x01,0x28,0x04,0x0f,0x57,0xfe,0x6c,0xfe,0x97,0x2a,0xb2,0x7d,0x84,0x10,0xc2,0x01,0x5c,0x34,0x06,0x11,0x9b,0x8c,0x2e,0xf6,0x05,0xc1,0x27,0xfd,0x21,0xfd,0x53,0x10,0x02,0x13,0x35,0x75,0x01,0x01,0x04,0x01,0x13,0x5f,0xfe,0xa1,0x0a,0x17,0x01,0x83,0x01,0x38,0xb2,0x72,0xfd,0xa6,0xd5,0x14,0x01,0x76,0x59,0x48,0x80,0x0b,0x46,0x00,0x00,0x00,0x02,0x00,0x9e,0xff,0xfe,0x01,0xa2,0x04,0x87,0x00,0x07,0x00,0x0f,0x00,0x00,0x36,0x37,0x32,0x17,0x14,0x07,0x26,0x27,0x12,0x37,0x32,0x17,0x14,0x07,0x26,0x27,0x9f,0x76,0x83,0x0a,0x7b,0x7f,0x0a,0x01,0x76,0x83,0x0a,0x7b,0x7f,0x0a,0xff,0x0a,0x7f,0x89,0x03,0x01,0x7a,0x04,0x04,0x0a,0x7f,0x89,0x03,0x01,0x7a,0x00,0x00,0x00,0x00,0x02,0x00,0x9e,0xff,0x08,0x01,0xa2,0x04,0x87,0x00,0x07,0x00,0x11,0x00,0x00,0x12,0x37,0x32,0x17,0x14,0x07,0x26,0x27,0x12,0x17,0x03,0x06,0x07,0x26,0x35,0x03,0x36,0x33,0x9f,0x76,0x83,0x0a,0x7b,0x7f,0x0a,0xdc,0x09,0x0d,0x01,0x57,0x57,0x0c,0x14,0x52,0x04,0x7d,0x0a,0x7f,0x89,0x03,0x01,0x7a,0xfc,0xfd,0x51,0xfe,0xd0,0x6a,0x01,0x01,0x6f,0x01,0x2f,0x51,0x00,0x00,0x00,0x01,0x00,0xc9,0x00,0x91,0x04,0x07,0x04,0x84,0x00,0x13,0x00,0x00,0x09,0x01,0x16,0x17,0x14,0x07,0x22,0x27,0x01,0x26,0x27,0x36,0x37,0x01,0x36,0x33,0x16,0x15,0x06,0x07,0x01,0xf6,0x01,0xc1,0x4e,0x02,0x46,0x3c,0x36,0xfd,0xd8,0x5b,0x03,0x03,0x5b,0x02,0x28,0x36,0x3c,0x46,0x02,0x4e,0x02,0x8b,0xfe,0xd6,0x27,0x4a,0x43,0x1c,0x20,0x01,0x56,0x1f,0x63,0x66,0x1f,0x01,0x56,0x20,0x1c,0x43,0x4a,0x27,0x00,0x00,0x00,0x02,0x00,0xc0,0x01,0x69,0x04,0x12,0x03,0x8b,0x00,0x09,0x00,0x13,0x00,0x00,0x00,0x17,0x06,0x07,0x05,0x26,0x27,0x36,0x33,0x25,0x12,0x17,0x06,0x07,0x21,0x26,0x27,0x36,0x33,0x25,0x04,0x04,0x0e,0x07,0x6c,0xfd,0x9b,0x75,0x05,0x08,0x73,0x02,0x5c,0x6d,0x0e,0x07,0x6c,0xfd,0x9b,0x75,0x05,0x08,0x73,0x02,0x5c,0x02,0x38,0x5e,0x62,0x0e,0x01,0x07,0x6b,0x5d,0x01,0x01,0x51,0x5f,0x62,0x0d,0x05,0x6b,0x5e,0x01,0x00,0x01,0x00,0xc9,0x00,0x91,0x04,0x07,0x04,0x84,0x00,0x13,0x00,0x00,0x01,0x26,0x27,0x34,0x37,0x32,0x17,0x01,0x16,0x17,0x06,0x07,0x01,0x06,0x23,0x26,0x35,0x36,0x37,0x01,0x01,0x19,0x4e,0x02,0x46,0x3c,0x36,0x02,0x28,0x5b,0x03,0x03,0x5b,0xfd,0xd8,0x36,0x3c,0x46,0x02,0x4e,0x01,0xc1,0x03,0xb4,0x27,0x4a,0x43,0x1c,0x20,0xfe,0xaa,0x1f,0x66,0x63,0x1f,0xfe,0xaa,0x20,0x1c,0x43,0x4a,0x27,0x01,0x2a,0x00,0x00,0x00,0x02,0x00,0xbc,0xff,0xff,0x03,0xca,0x07,0x4f,0x00,0x19,0x00,0x21,0x00,0x00,0x01,0x37,0x04,0x13,0x10,0x05,0x06,0x0f,0x01,0x06,0x23,0x26,0x35,0x34,0x37,0x36,0x35,0x34,0x27,0x0e,0x01,0x07,0x26,0x27,0x37,0x36,0x12,0x33,0x16,0x17,0x06,0x07,0x26,0x27,0x01,0xcf,0x79,0x01,0x74,0x0e,0xfe,0xb4,0x59,0x0a,0x01,0x15,0x61,0x63,0xbb,0xf9,0xe4,0x55,0x54,0x45,0x4c,0x1b,0x04,0x22,0x56,0x7b,0x63,0x1b,0x04,0x75,0x90,0x01,0x07,0x43,0x0c,0x14,0xfe,0x9a,0xfe,0xf5,0xe1,0x40,0x81,0xba,0x57,0x11,0xd7,0xf8,0x92,0x9e,0x9d,0xaa,0x09,0x0d,0x50,0x05,0x06,0x5d,0x2a,0x6b,0xfa,0x02,0x11,0x61,0x91,0x0d,0x19,0x8a,0x00,0x00,0x00,0x02,0x00,0x40,0x00,0x1e,0x06,0x10,0x05,0xa4,0x00,0x08,0x00,0x3d,0x00,0x00,0x01,0x14,0x17,0x36,0x13,0x27,0x37,0x06,0x08,0x01,0x05,0x26,0x2f,0x01,0x02,0x05,0x20,0x03,0x35,0x12,0x25,0x32,0x15,0x14,0x07,0x17,0x07,0x12,0x17,0x36,0x13,0x02,0x25,0x23,0x04,0x00,0x0f,0x01,0x12,0x05,0x36,0x37,0x17,0x16,0x17,0x16,0x17,0x06,0x07,0x26,0x27,0x05,0x24,0x03,0x27,0x12,0x00,0x25,0x37,0x04,0x13,0x17,0x01,0xcc,0x7e,0xe6,0xbd,0x04,0x04,0xe1,0xfe,0xd0,0x04,0x16,0xfe,0xfc,0xad,0x17,0x16,0xab,0xfe,0xf8,0xfe,0xe7,0x0b,0x3b,0x02,0x8c,0x91,0x0f,0x0f,0x02,0x09,0x56,0x7e,0x04,0x56,0xfe,0xf9,0x7e,0xfe,0xc9,0xfe,0x89,0x07,0x03,0x3a,0x01,0x3a,0xf1,0x77,0x66,0x95,0x98,0x2d,0x09,0x0e,0x54,0x8c,0x87,0xfe,0x43,0xfe,0x33,0x42,0x05,0x0d,0x01,0xd7,0x01,0x9b,0x4f,0x01,0x93,0x63,0x0c,0x02,0x64,0x94,0x16,0x05,0x01,0x54,0xc2,0x61,0x0b,0xfe,0xfc,0xfd,0xf8,0x08,0x0e,0xa9,0x82,0xfe,0xd4,0x04,0x01,0x20,0x47,0x02,0x1e,0x2b,0x4b,0x1f,0x17,0x81,0xcf,0xfe,0xb8,0x0b,0x38,0x01,0x50,0x01,0xd6,0x0c,0x10,0xfe,0x5c,0xd8,0x60,0xfe,0xb8,0x19,0x0a,0x05,0x04,0x07,0x16,0x0d,0x34,0x51,0x07,0x1e,0x0a,0x08,0x0d,0x01,0xb9,0x61,0x01,0x53,0x01,0xe0,0x0a,0x02,0x1c,0xfe,0x0a,0xa5,0x00,0x00,0x02,0x00,0x45,0xff,0xfc,0x06,0x62,0x07,0x4a,0x00,0x15,0x00,0x1c,0x00,0x00,0x01,0x04,0x00,0x13,0x11,0x14,0x23,0x22,0x35,0x11,0x21,0x11,0x14,0x07,0x26,0x27,0x11,0x36,0x37,0x16,0x15,0x12,0x03,0x21,0x26,0x00,0x21,0x20,0x00,0x03,0x81,0x01,0x77,0x01,0x67,0x03,0x5d,0x6e,0xfb,0x7d,0x67,0x67,0x01,0x04,0x60,0x6a,0xdc,0xbc,0x04,0x58,0x01,0xfe,0xff,0xfe,0xf3,0xfe,0xfb,0xfe,0xbc,0x07,0x4a,0x06,0xfe,0x13,0xfe,0x6a,0xfc,0x9f,0x64,0x62,0x02,0xff,0xfd,0x0d,0x6c,0x01,0x02,0x6b,0x05,0xb8,0x6c,0x01,0x01,0x90,0x01,0x4c,0xfc,0xd5,0xce,0x01,0x91,0xfe,0x64,0x00,0x00,0x00,0x00,0x02,0x00,0x57,0xff,0xf0,0x06,0x2f,0x07,0x65,0x00,0x25,0x00,0x2f,0x00,0x00,0x13,0x32,0x17,0x36,0x25,0x04,0x00,0x13,0x15,0x02,0x05,0x16,0x15,0x14,0x04,0x21,0x26,0x27,0x26,0x35,0x36,0x33,0x16,0x17,0x20,0x24,0x35,0x34,0x24,0x27,0x21,0x11,0x06,0x07,0x22,0x35,0x11,0x34,0x05,0x22,0x07,0x11,0x21,0x2c,0x01,0x37,0x26,0x00,0xb7,0x49,0x11,0x4e,0x01,0x01,0x01,0x81,0x02,0x3d,0x11,0x0b,0xfe,0xc3,0xcd,0xfe,0x5f,0xfe,0x6b,0x70,0x6d,0x55,0x02,0x65,0x65,0x6e,0x01,0x2a,0x01,0x3e,0xfe,0xe3,0xe4,0xfe,0x3b,0x21,0x51,0x5f,0x01,0xbf,0xe0,0x0e,0x01,0x75,0x01,0xa7,0x01,0x18,0x01,0x01,0xfe,0x2a,0x07,0x65,0x4d,0x2b,0x03,0x01,0xfe,0x74,0xfe,0xd0,0x31,0xfe,0xe3,0xb4,0x42,0xd8,0xc1,0xbc,0x07,0x08,0x1f,0x46,0x59,0x0c,0x02,0x63,0x62,0x67,0x48,0x03,0xfe,0x2a,0x50,0x0e,0x65,0x06,0xbc,0x4e,0xe3,0x2c,0xfc,0x9d,0x06,0xf4,0x9d,0xc4,0x01,0x33,0x00,0x01,0x00,0x3c,0xff,0xeb,0x05,0xe5,0x07,0x53,0x00,0x1a,0x00,0x00,0x01,0x32,0x04,0x17,0x06,0x07,0x22,0x26,0x23,0x06,0x00,0x03,0x12,0x00,0x33,0x20,0x36,0x33,0x16,0x17,0x14,0x04,0x05,0x24,0x03,0x12,0x00,0x03,0xb1,0xda,0x01,0x51,0x01,0x09,0x58,0x46,0xb7,0xd0,0xfa,0xfe,0x66,0x01,0x01,0x01,0x72,0xed,0x01,0x01,0xc2,0x52,0x55,0x01,0xfe,0x8d,0xff,0x00,0xfc,0xd0,0x06,0x02,0x02,0x18,0x07,0x53,0xbb,0x60,0x61,0x01,0x9d,0x01,0xfe,0x16,0xfe,0xbc,0xfe,0x9f,0xfe,0xe9,0x33,0x0f,0x5a,0x70,0x33,0x08,0x0d,0x03,0x55,0x01,0xbc,0x02,0x45,0x00,0x00,0x00,0x00,0x01,0x00,0x34,0xff,0xf2,0x06,0x11,0x07,0x65,0x00,0x1f,0x00,0x00,0x25,0x06,0x07,0x22,0x35,0x11,0x34,0x37,0x32,0x17,0x36,0x37,0x04,0x00,0x13,0x10,0x00,0x05,0x27,0x26,0x35,0x36,0x37,0x17,0x24,0x00,0x11,0x02,0x00,0x25,0x22,0x07,0x01,0x00,0x0d,0x5b,0x64,0x65,0x53,0x11,0x4e,0xf7,0x01,0x95,0x02,0x29,0x11,0xfd,0xf7,0xfe,0x62,0xfb,0x55,0x02,0x65,0xe7,0x01,0x43,0x01,0x94,0x01,0xfe,0x5c,0xfe,0x90,0xd6,0x54,0x50,0x50,0x0e,0x65,0x06,0xbc,0x4e,0x04,0x4d,0x2b,0x03,0x01,0xfe,0x74,0xfe,0x62,0xfe,0x81,0xfd,0x5f,0x02,0x06,0x1f,0x50,0x54,0x0a,0x05,0x15,0x01,0xf4,0x01,0x48,0x01,0x28,0x01,0x33,0x01,0x2c,0x00,0x00,0x01,0x00,0x38,0xff,0xfe,0x05,0x91,0x07,0x45,0x00,0x1a,0x00,0x00,0x01,0x16,0x15,0x06,0x07,0x21,0x03,0x21,0x16,0x15,0x06,0x07,0x21,0x11,0x21,0x16,0x15,0x06,0x07,0x21,0x26,0x27,0x11,0x26,0x27,0x34,0x37,0x04,0xef,0x5d,0x02,0x68,0xfc,0x47,0x01,0x03,0x5e,0x67,0x01,0x69,0xfc,0xa9,0x04,0x01,0x64,0x11,0x4e,0xfb,0x82,0x52,0x01,0x28,0x01,0x6a,0x07,0x45,0x09,0x58,0x66,0x03,0xfc,0x76,0x01,0x6b,0x5f,0x07,0xfe,0xa7,0x09,0x5b,0x57,0x0d,0x11,0x7f,0x05,0xf4,0x10,0x56,0x54,0x09,0x00,0x00,0x00,0x01,0x00,0x35,0xff,0xfd,0x04,0xa8,0x07,0x4c,0x00,0x16,0x00,0x00,0x01,0x16,0x15,0x06,0x07,0x21,0x11,0x21,0x16,0x15,0x06,0x07,0x21,0x13,0x06,0x07,0x26,0x27,0x11,0x26,0x27,0x34,0x37,0x04,0x4b,0x5d,0x02,0x68,0xfc,0xf0,0x02,0xa0,0x5d,0x01,0x5f,0xfd,0x65,0x01,0x06,0x69,0x63,0x01,0x28,0x01,0x6a,0x07,0x4c,0x09,0x58,0x68,0x03,0xfd,0x9d,0x0e,0x5f,0x61,0x07,0xfd,0x21,0x6b,0x01,0x01,0x72,0x06,0x19,0x10,0x56,0x54,0x09,0x00,0x00,0x01,0x00,0x1e,0xff,0xeb,0x07,0x19,0x07,0x53,0x00,0x28,0x00,0x00,0x01,0x13,0x21,0x22,0x27,0x36,0x37,0x21,0x16,0x17,0x14,0x07,0x27,0x11,0x06,0x23,0x26,0x2f,0x01,0x04,0x07,0x24,0x03,0x12,0x00,0x25,0x32,0x04,0x17,0x06,0x07,0x22,0x26,0x23,0x06,0x00,0x03,0x12,0x00,0x33,0x32,0x05,0x80,0x01,0xfe,0x9b,0x64,0x03,0x02,0x5f,0x02,0xae,0x53,0x02,0x51,0x7c,0x0f,0x5a,0x48,0x0f,0x03,0xfe,0xb7,0xf6,0xfc,0xda,0x06,0x02,0x02,0x18,0x01,0x5b,0xda,0x01,0x51,0x01,0x09,0x58,0x46,0xb7,0xd0,0xfa,0xfe,0x5c,0x01,0x01,0x01,0x68,0xf7,0xf7,0x01,0x81,0x01,0x0d,0x5d,0x66,0x03,0x0e,0x61,0x54,0x05,0x01,0xfd,0xb6,0x4b,0x04,0x44,0x4e,0x9b,0x08,0x0d,0x03,0x55,0x01,0xbc,0x02,0x45,0x05,0xbb,0x60,0x61,0x01,0x9d,0x01,0xfe,0x16,0xfe,0xbc,0xfe,0x9f,0xfe,0xe9,0x00,0x00,0x00,0x01,0x00,0x1d,0xff,0xf5,0x06,0xb7,0x07,0x47,0x00,0x22,0x00,0x00,0x01,0x13,0x36,0x37,0x32,0x17,0x11,0x16,0x15,0x06,0x07,0x11,0x06,0x23,0x26,0x27,0x03,0x21,0x11,0x06,0x23,0x26,0x27,0x11,0x26,0x35,0x36,0x37,0x11,0x36,0x37,0x32,0x17,0x11,0x21,0x05,0x8b,0x01,0x01,0x6d,0x6b,0x01,0x51,0x01,0x50,0x01,0x6b,0x6d,0x01,0x01,0xfb,0xc7,0x01,0x6b,0x6d,0x01,0x5b,0x02,0x59,0x01,0x6d,0x6b,0x01,0x04,0x39,0x03,0x6f,0x03,0x4d,0x8a,0x01,0x8a,0xfc,0x35,0x10,0x58,0x59,0x07,0xfe,0x50,0x85,0x01,0x85,0x01,0xab,0xfe,0x5a,0x81,0x01,0x81,0x01,0xaa,0x08,0x55,0x56,0x13,0x03,0xc8,0x8d,0x01,0x8c,0xfc,0x3b,0x00,0x00,0x00,0x00,0x01,0x00,0x33,0xff,0xfc,0x02,0x8f,0x07,0x44,0x00,0x17,0x00,0x00,0x13,0x23,0x22,0x35,0x34,0x33,0x21,0x32,0x15,0x14,0x2b,0x01,0x11,0x33,0x32,0x15,0x14,0x23,0x21,0x22,0x35,0x34,0x3b,0x01,0xf2,0x53,0x6c,0x71,0x01,0x7a,0x71,0x6c,0x5c,0x5c,0x6c,0x71,0xfe,0x86,0x71,0x6c,0x53,0x06,0x71,0x76,0x5d,0x5d,0x76,0xfa,0x5e,0x76,0x5d,0x5d,0x76,0x00,0x00,0x01,0x00,0x51,0xff,0xf6,0x06,0x9f,0x07,0x5b,0x00,0x21,0x00,0x00,0x01,0x05,0x26,0x35,0x36,0x33,0x21,0x34,0x37,0x32,0x17,0x33,0x32,0x15,0x06,0x2b,0x01,0x16,0x11,0x02,0x00,0x05,0x22,0x24,0x27,0x36,0x37,0x32,0x16,0x33,0x24,0x00,0x13,0x10,0x04,0xbb,0xfc,0x34,0x7f,0x06,0x78,0x03,0xa8,0x66,0x6e,0x01,0xb1,0x83,0x0a,0x6f,0x97,0x27,0x02,0xfe,0x42,0xfe,0x87,0xda,0xfe,0xaf,0x01,0x09,0x58,0x46,0xc2,0xd0,0x01,0x18,0x01,0x3f,0x01,0x06,0x10,0x01,0x01,0x69,0x6c,0x71,0x05,0x76,0x64,0x70,0xe4,0xfe,0xcf,0xfd,0xea,0xfe,0x15,0x05,0xbb,0x60,0x61,0x01,0xaa,0x01,0x01,0x89,0x01,0xb2,0x01,0x2c,0x00,0x01,0xff,0xf9,0xff,0xf8,0x06,0x46,0x07,0x53,0x00,0x24,0x00,0x00,0x01,0x00,0x01,0x36,0x37,0x16,0x15,0x14,0x07,0x00,0x01,0x04,0x01,0x16,0x15,0x06,0x07,0x26,0x27,0x00,0x25,0x11,0x14,0x23,0x22,0x27,0x33,0x03,0x26,0x27,0x34,0x37,0x03,0x34,0x33,0x32,0x15,0x01,0x1a,0x02,0xfe,0x01,0x64,0x1c,0x58,0x56,0x38,0xfe,0x7e,0xfc,0x98,0x02,0xf2,0x01,0xd6,0x4d,0x04,0x5f,0x3a,0x2f,0xfe,0x4c,0xfd,0x61,0x65,0x71,0x01,0x03,0x01,0x49,0x03,0x4c,0x01,0x71,0x65,0x03,0x5e,0x01,0x54,0x02,0x44,0x53,0x01,0x06,0x49,0x3f,0x61,0xfd,0x7d,0xfe,0xae,0x70,0xfe,0xc9,0x3f,0x52,0x4e,0x04,0x07,0x1d,0x01,0x27,0x6d,0xfe,0xa1,0x5d,0x5d,0x01,0xae,0x15,0x56,0x4f,0x25,0x04,0x07,0x6a,0x71,0x00,0x00,0x01,0x00,0x43,0xff,0xfa,0x05,0xa8,0x07,0x50,0x00,0x12,0x00,0x00,0x13,0x16,0x15,0x11,0x20,0x25,0x36,0x37,0x16,0x17,0x14,0x07,0x04,0x0d,0x01,0x26,0x27,0x03,0x36,0xaf,0x6d,0x02,0x7e,0x01,0x0f,0x4d,0x54,0x5a,0x04,0x7c,0xfe,0xe0,0xfe,0x9a,0xfe,0x67,0xc4,0x05,0x01,0x03,0x07,0x50,0x01,0x70,0xf9,0xf2,0x53,0x1f,0x0c,0x04,0x63,0x63,0x26,0x4c,0x16,0x03,0x09,0xbc,0x06,0x1d,0x73,0x00,0x00,0x01,0x00,0x3d,0x00,0x05,0x08,0xf0,0x07,0x43,0x00,0x1b,0x00,0x00,0x00,0x27,0x00,0x25,0x11,0x06,0x07,0x22,0x27,0x11,0x36,0x37,0x04,0x01,0x00,0x25,0x16,0x17,0x11,0x06,0x23,0x26,0x35,0x11,0x04,0x01,0x06,0x07,0x04,0x42,0x09,0xfe,0x99,0xfe,0x47,0x01,0x6d,0x61,0x0d,0x06,0x5d,0x02,0xb8,0x01,0x3f,0x01,0x3e,0x02,0xb8,0x5b,0x08,0x0d,0x61,0x70,0xfe,0x49,0xfe,0x99,0x09,0x56,0x01,0x2c,0x49,0x04,0x97,0x3d,0xfa,0x3f,0x82,0x01,0x86,0x06,0x45,0x6b,0x08,0x2f,0xfb,0xef,0x04,0x11,0x2f,0x08,0x6b,0xf9,0xbb,0x86,0x01,0x82,0x05,0xc1,0x3d,0xfb,0x69,0x49,0x05,0x00,0x00,0x00,0x00,0x01,0x00,0x3d,0xff,0xf7,0x06,0xc8,0x07,0x43,0x00,0x16,0x00,0x00,0x13,0x04,0x01,0x11,0x36,0x37,0x16,0x15,0x11,0x06,0x23,0x26,0x2f,0x01,0x00,0x25,0x11,0x14,0x07,0x22,0x27,0x11,0x36,0xa0,0x03,0xa3,0x01,0xaa,0x02,0x5b,0x7e,0x08,0x63,0x62,0x09,0x01,0xfe,0x35,0xfc,0xf0,0x6b,0x61,0x0d,0x06,0x07,0x43,0x57,0xfc,0x47,0x03,0x91,0x60,0x18,0x01,0x79,0xf9,0x9e,0x69,0x0a,0x57,0xcd,0x04,0xbf,0x6f,0xfa,0x35,0x82,0x01,0x86,0x06,0x45,0x6b,0x00,0x00,0x00,0x02,0x00,0x1a,0xff,0xe4,0x07,0x7f,0x07,0x5a,0x00,0x13,0x00,0x25,0x00,0x00,0x01,0x16,0x17,0x06,0x23,0x22,0x26,0x27,0x22,0x00,0x03,0x12,0x00,0x05,0x20,0x00,0x13,0x10,0x00,0x2d,0x01,0x26,0x35,0x34,0x37,0x36,0x37,0x04,0x00,0x13,0x02,0x00,0x21,0x24,0x00,0x11,0x12,0x00,0x03,0x3d,0xc1,0x01,0x0a,0x51,0x31,0x6e,0x6c,0x77,0xfe,0xd9,0x02,0x0a,0x01,0xa7,0x01,0x0f,0x01,0x0c,0x01,0xc0,0x15,0xfe,0x35,0xfe,0xe7,0xfe,0x56,0x27,0x3c,0xaa,0xed,0x01,0x84,0x02,0x42,0x01,0x23,0xfd,0xfa,0xfe,0x62,0xfe,0x70,0xfd,0xf2,0x02,0x01,0x6d,0x06,0x92,0x22,0x7d,0x3f,0x50,0x01,0xfe,0x7b,0xfe,0xf5,0xfe,0x81,0xfe,0xc0,0x05,0x01,0x2c,0x01,0x94,0x01,0xb3,0x01,0x71,0x09,0x08,0x0b,0x43,0x25,0x24,0x15,0x08,0x09,0xfe,0x33,0xfd,0xe8,0xfe,0x2c,0xfe,0x4c,0x01,0x01,0xe8,0x01,0xaa,0x01,0x40,0x01,0xef,0x00,0x00,0x00,0x02,0x00,0x3d,0xff,0xf2,0x06,0x25,0x07,0x65,0x00,0x13,0x00,0x1d,0x00,0x00,0x00,0x29,0x01,0x11,0x06,0x07,0x22,0x35,0x11,0x34,0x37,0x32,0x17,0x36,0x25,0x04,0x00,0x13,0x15,0x06,0x01,0x22,0x07,0x11,0x21,0x24,0x36,0x37,0x26,0x00,0x04,0x7a,0xfe,0x69,0xfe,0x27,0x0d,0x5c,0x64,0x65,0x54,0x11,0x4e,0x01,0x01,0x01,0x95,0x02,0x29,0x11,0x0b,0xfc,0x24,0xe0,0x54,0x01,0xbb,0x01,0x9d,0xf0,0x01,0x01,0xfe,0x5c,0x02,0x22,0xfe,0x2e,0x50,0x0e,0x65,0x06,0xbc,0x4e,0x04,0x4d,0x2b,0x03,0x01,0xfe,0x74,0xfe,0xd0,0x31,0xff,0x03,0x1b,0x2c,0xfc,0xa7,0x06,0xea,0x9d,0xc4,0x01,0x33,0x00,0x02,0x00,0x24,0xfe,0x33,0x07,0xa6,0x07,0x5a,0x00,0x16,0x00,0x2e,0x00,0x00,0x25,0x26,0x27,0x36,0x33,0x16,0x17,0x16,0x33,0x32,0x00,0x13,0x02,0x00,0x25,0x20,0x00,0x03,0x10,0x00,0x05,0x37,0x26,0x04,0x05,0x16,0x17,0x06,0x07,0x26,0x27,0x26,0x27,0x06,0x07,0x24,0x00,0x03,0x12,0x00,0x21,0x04,0x00,0x11,0x02,0x00,0x07,0x03,0xc4,0x33,0x03,0x04,0x68,0x51,0x34,0x61,0x20,0x77,0x01,0x27,0x02,0x0a,0xfe,0x59,0xfe,0xf1,0xfe,0xf4,0xfe,0x40,0x15,0x01,0xcb,0x01,0x19,0x56,0x3e,0x02,0x53,0x01,0x07,0x4d,0x04,0x11,0x4c,0x5b,0x57,0xe9,0x9a,0x88,0xab,0xfe,0x68,0xfd,0xdc,0x01,0x23,0x01,0xfc,0x01,0x9e,0x01,0x90,0x02,0x04,0x02,0xfe,0xa7,0x83,0xeb,0x21,0x44,0x58,0x02,0x37,0x36,0x01,0x86,0x01,0x0a,0x01,0x7f,0x01,0x40,0x05,0xfe,0xd4,0xfe,0x6c,0xfe,0x4d,0xfe,0x8f,0x08,0x08,0x1d,0xdc,0xde,0x3b,0x42,0x4f,0x0d,0x02,0x67,0xd3,0x87,0x16,0x06,0x09,0x01,0xe2,0x02,0x0d,0x01,0xd4,0x01,0xb4,0x01,0xfe,0x18,0xfe,0x56,0xfe,0xb6,0xfe,0x1b,0x14,0x00,0x00,0x02,0x00,0x27,0xff,0xf2,0x06,0x3b,0x07,0x65,0x00,0x19,0x00,0x22,0x00,0x00,0x13,0x32,0x17,0x36,0x25,0x04,0x00,0x13,0x02,0x05,0x01,0x16,0x15,0x14,0x23,0x26,0x27,0x01,0x21,0x11,0x06,0x07,0x22,0x35,0x11,0x34,0x05,0x22,0x07,0x11,0x21,0x20,0x13,0x26,0x00,0x96,0x4c,0x11,0x4e,0x01,0x01,0x01,0x95,0x02,0x29,0x11,0x01,0xfe,0x9c,0x01,0x71,0x1e,0x70,0x57,0x42,0xfe,0x8b,0xfd,0x39,0x0d,0x54,0x6e,0x02,0x03,0xe0,0x54,0x02,0x01,0x02,0x3d,0x01,0x01,0xfe,0x66,0x07,0x65,0x4d,0x2b,0x03,0x01,0xfe,0x74,0xfe,0xd0,0xfe,0x6c,0x90,0xfe,0x3f,0x26,0x2c,0x5c,0x01,0x70,0x01,0xbf,0xfe,0x2a,0x50,0x0e,0x65,0x06,0xbc,0x4e,0xf4,0x25,0xfc,0xa7,0x01,0x8d,0xc4,0x01,0x2c,0x00,0x00,0x00,0x00,0x01,0x00,0x2a,0xff,0xe3,0x06,0x0b,0x07,0x5c,0x00,0x21,0x00,0x00,0x01,0x04,0x17,0x16,0x17,0x06,0x07,0x22,0x26,0x25,0x04,0x03,0x16,0x00,0x13,0x02,0x05,0x24,0x27,0x26,0x27,0x36,0x37,0x32,0x17,0x16,0x05,0x24,0x37,0x34,0x24,0x03,0x12,0x25,0x03,0x63,0x01,0x70,0xe5,0x52,0x01,0x10,0x46,0x3f,0xcc,0xfe,0xb5,0xfd,0xa8,0x07,0x01,0x04,0xd9,0x01,0x16,0xfd,0x89,0xfe,0x6e,0xd8,0x52,0x01,0x06,0x50,0x2b,0x4e,0xcc,0x01,0x26,0x01,0xa3,0x0b,0xfb,0x2b,0x01,0x1a,0x03,0x1e,0x07,0x5c,0x02,0x91,0x34,0x53,0x57,0x01,0xa0,0x0b,0x1f,0xfe,0x73,0xf4,0xfe,0xf9,0xfe,0x8c,0xfe,0x7d,0x14,0x11,0x85,0x3e,0x44,0x66,0x01,0x3f,0x6a,0x07,0x1d,0xaf,0xe5,0xf4,0x01,0x97,0x02,0x54,0x1a,0x00,0x00,0x01,0x00,0x01,0xff,0xfc,0x05,0x91,0x07,0x44,0x00,0x10,0x00,0x00,0x01,0x21,0x22,0x35,0x34,0x33,0x21,0x32,0x15,0x14,0x23,0x21,0x03,0x14,0x23,0x22,0x27,0x02,0x61,0xfe,0x0c,0x6c,0x71,0x04,0xae,0x71,0x6c,0xfe,0x17,0x02,0x67,0x71,0x01,0x06,0x71,0x76,0x5d,0x5d,0x76,0xf9,0xe8,0x5d,0x5d,0x00,0x00,0x00,0x00,0x01,0x00,0x16,0xff,0xfc,0x06,0x02,0x07,0x5b,0x00,0x1b,0x00,0x00,0x13,0x36,0x33,0x16,0x17,0x02,0x11,0x12,0x00,0x05,0x32,0x37,0x11,0x36,0x33,0x32,0x15,0x11,0x14,0x07,0x22,0x27,0x06,0x07,0x24,0x00,0x03,0x10,0x63,0x0c,0x64,0x68,0x01,0x4a,0x01,0x01,0x9a,0x01,0x70,0xcc,0x5e,0x0d,0x64,0x6a,0x65,0x62,0x11,0x58,0xed,0xfe,0x6b,0xfd,0xd7,0x11,0x06,0xdf,0x74,0x02,0x79,0xfd,0x7d,0xfe,0xd6,0xfe,0xd8,0xfe,0xcd,0x01,0x54,0x05,0xcb,0x6d,0x6f,0xf9,0x62,0x4e,0x04,0x4d,0x49,0x03,0x01,0x01,0x8c,0x01,0x9e,0x01,0x48,0x00,0x00,0x00,0x00,0x01,0x00,0x02,0xff,0xfe,0x06,0x43,0x07,0x48,0x00,0x14,0x00,0x00,0x09,0x01,0x36,0x33,0x16,0x15,0x06,0x07,0x01,0x06,0x07,0x23,0x26,0x27,0x01,0x26,0x27,0x34,0x37,0x32,0x17,0x03,0x23,0x02,0x3b,0x2a,0x5a,0x61,0x08,0x18,0xfd,0x85,0x26,0x5f,0x01,0x5f,0x26,0xfd,0x85,0x18,0x08,0x57,0x64,0x2a,0x01,0x64,0x05,0x60,0x84,0x10,0x69,0x37,0x35,0xfa,0x14,0x76,0x03,0x03,0x76,0x05,0xec,0x35,0x37,0x69,0x10,0x84,0x00,0x01,0x00,0x02,0xff,0xfe,0x09,0x63,0x07,0x48,0x00,0x29,0x00,0x00,0x09,0x01,0x06,0x07,0x23,0x26,0x27,0x01,0x26,0x27,0x34,0x37,0x32,0x17,0x09,0x01,0x36,0x37,0x36,0x37,0x32,0x17,0x36,0x33,0x16,0x17,0x16,0x17,0x09,0x01,0x36,0x33,0x16,0x15,0x06,0x07,0x01,0x06,0x07,0x23,0x26,0x27,0x04,0xb3,0xfe,0xf5,0x26,0x5f,0x01,0x5f,0x26,0xfd,0x85,0x18,0x08,0x57,0x67,0x2a,0x02,0x39,0x01,0x19,0x0a,0x0d,0x10,0x42,0x07,0x06,0x07,0x07,0x42,0x10,0x0d,0x0a,0x01,0x1a,0x02,0x37,0x2a,0x64,0x5b,0x08,0x18,0xfd,0x85,0x26,0x5f,0x01,0x5f,0x26,0x02,0xd0,0xfd,0xa7,0x76,0x03,0x03,0x76,0x05,0xec,0x35,0x37,0x69,0x10,0x84,0xfa,0xa0,0x02,0x68,0x20,0x18,0x40,0x0c,0x01,0x01,0x0c,0x40,0x18,0x20,0xfd,0x98,0x05,0x60,0x84,0x10,0x69,0x37,0x35,0xfa,0x14,0x76,0x03,0x03,0x76,0x00,0x01,0x00,0x12,0xff,0xf4,0x05,0x53,0x07,0x4f,0x00,0x1f,0x00,0x00,0x09,0x01,0x26,0x27,0x34,0x37,0x32,0x17,0x09,0x01,0x36,0x33,0x16,0x15,0x06,0x07,0x09,0x01,0x16,0x17,0x14,0x07,0x22,0x27,0x09,0x01,0x06,0x23,0x26,0x35,0x36,0x37,0x01,0xf9,0xfe,0x40,0x1d,0x0a,0x53,0x63,0x37,0x01,0xaf,0x01,0xb8,0x37,0x63,0x53,0x0a,0x1d,0xfe,0x37,0x01,0xc9,0x1d,0x0a,0x53,0x63,0x37,0xfe,0x48,0xfe,0x51,0x37,0x63,0x53,0x0a,0x1d,0x03,0xa2,0x02,0xc8,0x35,0x37,0x69,0x10,0x84,0xfd,0x5f,0x02,0x97,0x84,0x10,0x69,0x37,0x35,0xfd,0x42,0xfd,0x41,0x35,0x37,0x69,0x10,0x84,0x02,0x97,0xfd,0x5f,0x84,0x10,0x69,0x37,0x35,0x00,0x00,0x00,0x01,0x00,0x21,0xff,0xff,0x05,0xc0,0x07,0x4f,0x00,0x15,0x00,0x00,0x09,0x01,0x26,0x27,0x34,0x37,0x32,0x17,0x09,0x01,0x36,0x33,0x16,0x15,0x06,0x07,0x01,0x11,0x14,0x07,0x26,0x27,0x02,0x7d,0xfd,0xcd,0x1f,0x0a,0x64,0x5f,0x36,0x01,0xd2,0x01,0xdb,0x36,0x5f,0x64,0x0a,0x1f,0xfd,0xc2,0x6d,0x6e,0x01,0x02,0x23,0x04,0x47,0x35,0x37,0x69,0x10,0x84,0xfc,0x76,0x03,0x80,0x84,0x10,0x69,0x37,0x35,0xfb,0xc3,0xfe,0x4d,0x6a,0x07,0x07,0x6a,0x00,0x00,0x00,0x00,0x01,0x00,0x31,0xff,0xfe,0x05,0xb9,0x07,0x3f,0x00,0x17,0x00,0x00,0x08,0x01,0x35,0x21,0x22,0x27,0x36,0x37,0x25,0x16,0x15,0x02,0x00,0x06,0x15,0x05,0x32,0x17,0x06,0x07,0x21,0x26,0x35,0x10,0x01,0x43,0x03,0x83,0xfb,0xf9,0x7f,0x0f,0x06,0x88,0x04,0x7a,0x80,0x0a,0xfc,0x5a,0xdb,0x03,0xdf,0x7f,0x0f,0x06,0x88,0xfb,0xa4,0x80,0x02,0xb8,0x02,0xb5,0xfc,0x67,0x69,0x05,0x01,0x0b,0x87,0xfe,0x7a,0xfd,0x17,0xe7,0x7a,0x01,0x71,0x68,0x05,0x09,0x87,0x01,0x02,0x00,0x00,0x00,0x00,0x01,0x00,0xaa,0xff,0x21,0x02,0xd0,0x08,0x26,0x00,0x11,0x00,0x00,0x13,0x34,0x33,0x25,0x16,0x15,0x06,0x07,0x21,0x11,0x25,0x16,0x17,0x14,0x07,0x25,0x22,0x35,0xaa,0x6c,0x01,0x50,0x6a,0x02,0x5c,0xfe,0xec,0x01,0x14,0x5c,0x02,0x6a,0xfe,0xb0,0x6c,0x07,0xa1,0x83,0x02,0x0b,0x4e,0x67,0x02,0xf8,0x7f,0x01,0x02,0x68,0x4e,0x0b,0x02,0x83,0x00,0x00,0x00,0x01,0x00,0x0f,0xff,0x8e,0x03,0x07,0x07,0xf9,0x00,0x0d,0x00,0x00,0x12,0x37,0x16,0x17,0x01,0x16,0x15,0x06,0x07,0x26,0x27,0x01,0x26,0x35,0x0f,0x6c,0x4f,0x0c,0x02,0x1a,0x17,0x0b,0x46,0x48,0x1a,0xfd,0xe1,0x26,0x07,0xf7,0x02,0x11,0x5e,0xf8,0xcb,0x2a,0x44,0x58,0x01,0x05,0x42,0x07,0x32,0x41,0x54,0x00,0x00,0x01,0x00,0x50,0xff,0x21,0x02,0x76,0x08,0x26,0x00,0x11,0x00,0x00,0x05,0x14,0x23,0x05,0x26,0x35,0x36,0x37,0x05,0x11,0x21,0x26,0x27,0x34,0x37,0x05,0x32,0x15,0x02,0x76,0x6c,0xfe,0xb0,0x6a,0x02,0x5c,0x01,0x14,0xfe,0xec,0x5c,0x02,0x6a,0x01,0x50,0x6c,0x5a,0x83,0x02,0x0b,0x4e,0x68,0x02,0x01,0x07,0x81,0x02,0x67,0x4e,0x0b,0x02,0x83,0x00,0x00,0x00,0x01,0xff,0xa6,0xfe,0xdd,0x04,0xd8,0xff,0x90,0x00,0x09,0x00,0x00,0x01,0x21,0x26,0x27,0x36,0x33,0x21,0x32,0x15,0x06,0x04,0x76,0xfb,0x90,0x5e,0x02,0x02,0x5d,0x04,0x72,0x61,0x02,0xfe,0xdd,0x01,0x5d,0x55,0x5c,0x56,0x00,0x00,0x01,0x00,0x4a,0x05,0x23,0x02,0x6b,0x06,0x13,0x00,0x0e,0x00,0x00,0x00,0x15,0x06,0x07,0x26,0x25,0x26,0x27,0x36,0x33,0x32,0x17,0x1e,0x01,0x17,0x02,0x6b,0x01,0x34,0x87,0xfe,0xd5,0x37,0x03,0x07,0x3e,0x34,0x4b,0xa9,0x62,0x21,0x05,0x82,0x2a,0x2d,0x08,0x07,0x6c,0x16,0x2a,0x3d,0x2a,0x3b,0x0f,0x0b,0x00,0x00,0x02,0x00,0x3e,0xff,0xf9,0x04,0xca,0x04,0x93,0x00,0x09,0x00,0x26,0x00,0x00,0x25,0x36,0x24,0x37,0x34,0x25,0x06,0x04,0x07,0x16,0x01,0x13,0x06,0x07,0x26,0x2f,0x01,0x06,0x21,0x24,0x03,0x36,0x00,0x25,0x32,0x17,0x2e,0x01,0x27,0x22,0x06,0x23,0x26,0x35,0x36,0x24,0x37,0x04,0x12,0x01,0xb0,0xc0,0x01,0x6c,0x07,0xfe,0xf3,0xaa,0xfe,0xd8,0x01,0x06,0x03,0xad,0x14,0x07,0x5f,0x55,0x0a,0x06,0xef,0xfe,0x8b,0xfe,0xa6,0x03,0x01,0x01,0x8c,0x01,0x00,0xd2,0x4e,0x01,0x83,0xb7,0xcd,0x8e,0x4d,0x49,0x06,0x01,0x15,0xdb,0x01,0x27,0xd9,0xb9,0x0c,0x98,0x80,0x7d,0x0a,0x06,0xaa,0x6e,0x8d,0x02,0x0c,0xfd,0xb5,0x70,0x0a,0x09,0x40,0x63,0xb3,0x12,0x01,0x39,0xb6,0x01,0x10,0x14,0x2d,0x5d,0x77,0x0c,0x69,0x08,0x60,0x4e,0x70,0x05,0x07,0xfe,0xf5,0x00,0x00,0x02,0x00,0x4b,0xff,0xef,0x04,0xce,0x07,0x56,0x00,0x09,0x00,0x1c,0x00,0x00,0x01,0x06,0x00,0x07,0x14,0x33,0x36,0x00,0x37,0x26,0x01,0x36,0x37,0x16,0x17,0x11,0x12,0x21,0x04,0x13,0x02,0x00,0x05,0x22,0x27,0x06,0x23,0x22,0x27,0x03,0x5c,0xc0,0xfe,0x94,0x07,0xd8,0xad,0x01,0x3f,0x17,0x06,0xfc,0x4d,0x03,0x67,0x61,0x01,0xe5,0x01,0x6b,0x01,0x5a,0x0d,0x01,0xfe,0x74,0xfe,0xc4,0x96,0x58,0x1e,0x56,0x57,0x01,0x03,0x9e,0x02,0xfe,0x82,0x9e,0xcd,0x01,0x01,0x31,0xf0,0xc9,0x03,0x44,0x73,0x01,0x02,0x80,0xfc,0x37,0x01,0x5d,0x12,0xfe,0x81,0xfe,0xf8,0xfe,0x34,0x14,0x26,0x26,0x71,0x00,0x00,0x00,0x00,0x01,0x00,0x39,0xff,0xec,0x04,0x10,0x04,0x88,0x00,0x19,0x00,0x00,0x01,0x04,0x17,0x06,0x07,0x2e,0x01,0x23,0x0e,0x01,0x07,0x12,0x17,0x3e,0x02,0x37,0x16,0x17,0x06,0x04,0x07,0x24,0x03,0x12,0x00,0x02,0x6c,0x01,0x64,0x05,0x02,0x58,0x35,0x7d,0x58,0x83,0xee,0x02,0x14,0xf4,0x8d,0xb8,0x2b,0x47,0x4d,0x06,0x09,0xfe,0xeb,0xdd,0xfe,0x2f,0x0b,0x01,0x01,0x1e,0x04,0x88,0x0b,0x99,0x53,0x05,0x01,0x37,0x01,0xff,0xbf,0xfe,0xb5,0x06,0x01,0xa5,0x63,0x01,0x04,0x64,0x74,0xf1,0x05,0x05,0x01,0xfc,0x01,0x1f,0x01,0x67,0x00,0x02,0x00,0x34,0xff,0xf9,0x04,0xe8,0x07,0x47,0x00,0x0a,0x00,0x20,0x00,0x00,0x25,0x36,0x00,0x37,0x27,0x34,0x23,0x06,0x00,0x07,0x16,0x01,0x03,0x36,0x37,0x16,0x17,0x1a,0x01,0x17,0x06,0x07,0x26,0x35,0x27,0x02,0x21,0x24,0x03,0x12,0x00,0x25,0x32,0x01,0xa6,0xc0,0x01,0x6c,0x0a,0x03,0xd8,0xad,0xfe,0xc1,0x1c,0x06,0x02,0xe5,0x06,0x03,0x6f,0x5a,0x05,0x05,0x33,0x01,0x07,0x5f,0x69,0x1a,0xf9,0xfe,0x8b,0xfe,0xa6,0x03,0x01,0x01,0x8c,0x01,0x3c,0x90,0xb9,0x0c,0x01,0x7e,0x98,0x56,0x7d,0x01,0xfe,0xcf,0xf0,0xd3,0x03,0x96,0x02,0x80,0x76,0x02,0x0e,0x6b,0xfc,0x91,0xfd,0x76,0x5b,0x70,0x0a,0x09,0x72,0xf9,0xfe,0x85,0x12,0x01,0x7f,0x01,0x08,0x01,0xcc,0x14,0x00,0x02,0x00,0x39,0xff,0xec,0x04,0x82,0x04,0x93,0x00,0x07,0x00,0x1d,0x00,0x00,0x01,0x34,0x23,0x04,0x07,0x16,0x17,0x20,0x16,0x05,0x26,0x27,0x12,0x05,0x36,0x37,0x36,0x33,0x16,0x17,0x06,0x04,0x05,0x24,0x03,0x12,0x00,0x25,0x04,0x13,0x03,0xb3,0xd7,0xfe,0xba,0x57,0x93,0x66,0x01,0x78,0xcb,0xfd,0xc7,0xbf,0x6c,0x09,0x01,0x64,0xa0,0x88,0x41,0x41,0x53,0x01,0x02,0xfe,0xdd,0xfe,0xdc,0xfe,0x27,0x27,0x01,0x01,0x7e,0x01,0x23,0x01,0x9d,0x04,0x03,0x4c,0x88,0x1c,0xd4,0x08,0x02,0xbc,0x0c,0x0a,0x01,0xfe,0xaa,0x13,0x02,0x78,0x3d,0x01,0x60,0x4e,0xce,0x02,0x38,0x01,0xe0,0x01,0x27,0x01,0x5b,0x0d,0x0f,0xfe,0xcc,0x00,0x00,0x01,0xff,0xc6,0x00,0x00,0x02,0x9d,0x07,0x49,0x00,0x1e,0x00,0x00,0x01,0x1e,0x01,0x17,0x06,0x07,0x2e,0x01,0x27,0x06,0x07,0x33,0x16,0x17,0x06,0x07,0x23,0x13,0x14,0x07,0x22,0x27,0x03,0x23,0x22,0x35,0x34,0x3f,0x01,0x3e,0x01,0x01,0x8c,0x87,0x89,0x01,0x08,0x46,0x1e,0x60,0x4a,0x64,0x04,0xeb,0x4d,0x04,0x08,0x4d,0xea,0x0b,0x64,0x60,0x0e,0x0d,0x2d,0x55,0x5a,0x31,0x05,0x94,0x07,0x49,0x01,0x48,0x47,0x4a,0x02,0x01,0x1b,0x02,0x0c,0xce,0x0b,0x42,0x5a,0x08,0xfb,0x79,0x70,0x0b,0x7c,0x04,0x85,0x5b,0x4f,0x05,0x04,0xac,0xe8,0x00,0x00,0x02,0x00,0x27,0xfd,0xe4,0x04,0xbf,0x04,0x68,0x00,0x0a,0x00,0x28,0x00,0x00,0x25,0x36,0x00,0x37,0x27,0x34,0x23,0x06,0x00,0x07,0x16,0x08,0x01,0x07,0x2e,0x01,0x35,0x36,0x37,0x32,0x16,0x33,0x3e,0x01,0x37,0x13,0x02,0x21,0x24,0x03,0x12,0x00,0x25,0x32,0x17,0x36,0x33,0x16,0x17,0x13,0x03,0x01,0x99,0xc0,0x01,0x6c,0x0a,0x03,0xd8,0xad,0xfe,0xc1,0x1c,0x06,0x03,0xc4,0xfe,0xd7,0xe7,0xc0,0xa9,0x03,0x56,0x4f,0x6d,0x59,0x67,0xde,0x02,0x03,0xfc,0xfe,0x8b,0xfe,0xa6,0x03,0x01,0x01,0x8c,0x01,0x3c,0x96,0x58,0x1e,0x55,0x61,0x01,0x0c,0x09,0xaf,0x0c,0x01,0x7e,0x98,0x56,0x7d,0x01,0xfe,0xcf,0xf0,0xd3,0xfe,0x82,0xfe,0xb8,0x05,0x01,0x4d,0x50,0x45,0x14,0x30,0x01,0xc3,0xe9,0x01,0x12,0xfe,0x85,0x12,0x01,0x7f,0x01,0x08,0x01,0xcc,0x14,0x26,0x26,0x01,0x70,0xfd,0xeb,0xfe,0x58,0x00,0x00,0x01,0x00,0x42,0x00,0x03,0x04,0x66,0x07,0x3d,0x00,0x1b,0x00,0x00,0x37,0x26,0x35,0x02,0x35,0x36,0x37,0x16,0x17,0x13,0x12,0x25,0x04,0x13,0x14,0x03,0x06,0x23,0x26,0x35,0x12,0x35,0x26,0x27,0x22,0x00,0x03,0x06,0xc5,0x67,0x1c,0x0d,0x58,0x60,0x07,0x09,0x9e,0x01,0x4f,0x01,0x5d,0x05,0x14,0x0a,0x68,0x55,0x10,0x0a,0x93,0x92,0xfe,0xf4,0x32,0x05,0x07,0x0c,0x68,0x06,0x17,0x4c,0x5e,0x01,0x09,0x7a,0xfc,0x5a,0x01,0x6d,0x07,0x0a,0xfe,0x44,0xf2,0xfe,0x98,0x65,0x08,0x63,0x01,0x66,0xdf,0xfd,0x11,0xfe,0x83,0xfe,0x2a,0x5e,0x00,0x00,0x00,0x02,0x00,0x52,0xff,0xf9,0x02,0x3e,0x06,0x99,0x00,0x07,0x00,0x18,0x00,0x00,0x01,0x16,0x15,0x06,0x07,0x26,0x27,0x36,0x12,0x17,0x03,0x16,0x33,0x32,0x36,0x33,0x32,0x17,0x06,0x07,0x24,0x03,0x13,0x36,0x33,0x01,0x05,0x69,0x13,0x65,0x72,0x02,0x16,0x8d,0x01,0x09,0x14,0x5d,0x1c,0x33,0x22,0x35,0x0a,0x02,0xbc,0xfe,0xd7,0x05,0x0b,0x05,0x62,0x06,0x99,0x1a,0x6c,0x68,0x0c,0x05,0x8f,0x66,0xfd,0xe5,0x6d,0xfd,0x8f,0xda,0x12,0x4f,0x8f,0x01,0x17,0x01,0x9a,0x02,0x69,0x6b,0x00,0x02,0xfe,0xb5,0xfe,0x5c,0x01,0x9c,0x07,0x12,0x00,0x08,0x00,0x1b,0x00,0x00,0x01,0x16,0x17,0x07,0x06,0x23,0x22,0x27,0x34,0x13,0x16,0x17,0x13,0x0a,0x01,0x07,0x24,0x27,0x36,0x37,0x32,0x16,0x33,0x32,0x36,0x13,0x03,0x36,0x01,0x06,0x80,0x0a,0x0a,0x27,0x58,0x5b,0x13,0x8a,0x4f,0x13,0x17,0x01,0xe3,0xf2,0xff,0x00,0x11,0x03,0x3d,0x2e,0x56,0x51,0x82,0x84,0x01,0x15,0x05,0x07,0x12,0x01,0x6c,0x3d,0x5d,0x70,0x7d,0xfd,0x9d,0x03,0x69,0xfc,0xed,0xfe,0x78,0xfe,0xd4,0x06,0x10,0x85,0x54,0x0c,0x26,0xca,0x01,0x41,0x02,0xfa,0x57,0x00,0x00,0x01,0x00,0x3e,0xff,0xf9,0x04,0x2e,0x07,0x2b,0x00,0x1b,0x00,0x00,0x12,0x37,0x32,0x15,0x03,0x01,0x36,0x37,0x32,0x17,0x06,0x07,0x05,0x01,0x16,0x17,0x06,0x07,0x26,0x27,0x01,0x07,0x13,0x06,0x23,0x26,0x27,0x13,0x4b,0x6f,0x66,0x09,0x01,0xda,0x50,0x3b,0x68,0x07,0x08,0x7c,0xfe,0xcf,0x01,0xd9,0x1e,0x01,0x03,0x52,0x57,0x15,0xfe,0x0e,0x5b,0x02,0x01,0x6b,0x75,0x03,0x0b,0x07,0x23,0x08,0x6f,0xfc,0x3f,0x01,0x31,0x43,0x01,0x73,0x45,0x3d,0xc5,0xfd,0xfb,0x24,0x3f,0x4a,0x0b,0x0b,0x2a,0x02,0x21,0x3d,0xfe,0x6f,0x81,0x01,0x78,0x06,0x32,0x00,0x00,0x00,0x00,0x01,0x00,0x38,0xff,0xf9,0x02,0x24,0x07,0x4a,0x00,0x10,0x00,0x00,0x00,0x17,0x03,0x16,0x33,0x32,0x36,0x33,0x32,0x17,0x06,0x07,0x24,0x03,0x13,0x36,0x33,0x01,0x10,0x01,0x0e,0x14,0x5d,0x1c,0x33,0x22,0x35,0x0a,0x02,0xbc,0xfe,0xd7,0x05,0x10,0x05,0x62,0x07,0x4a,0x6d,0xfa,0xc3,0xda,0x12,0x4f,0x8f,0x01,0x17,0x01,0x9a,0x05,0x35,0x6b,0x00,0x00,0x00,0x01,0x00,0x46,0xff,0xfa,0x07,0x41,0x04,0x88,0x00,0x2e,0x00,0x00,0x01,0x06,0x03,0x06,0x23,0x26,0x35,0x12,0x35,0x26,0x27,0x22,0x00,0x03,0x06,0x07,0x26,0x35,0x0a,0x01,0x35,0x36,0x37,0x16,0x17,0x13,0x12,0x25,0x16,0x17,0x36,0x37,0x04,0x13,0x14,0x03,0x06,0x23,0x26,0x35,0x12,0x35,0x26,0x27,0x22,0x07,0x06,0x04,0x85,0x03,0x11,0x0a,0x68,0x55,0x10,0x0a,0x93,0x92,0xfe,0xf4,0x32,0x05,0x66,0x67,0x07,0x2e,0x0d,0x58,0x6a,0x07,0x10,0xa8,0x01,0x4f,0xe5,0x51,0x99,0xed,0x01,0x5d,0x05,0x14,0x0a,0x68,0x55,0x10,0x0a,0x93,0x92,0x86,0x21,0x02,0x92,0xe6,0xfe,0xb9,0x65,0x08,0x63,0x01,0x66,0xdf,0xfd,0x11,0xfe,0x83,0xfe,0x20,0x5e,0x09,0x0c,0x68,0x01,0xcd,0x01,0xa2,0x4c,0x5e,0x01,0x09,0x7a,0xfe,0xf8,0x01,0x81,0x07,0x07,0xc0,0xc2,0x05,0x0a,0xfe,0x44,0xf2,0xfe,0x98,0x65,0x08,0x63,0x01,0x66,0xdf,0xfd,0x11,0xbe,0x2f,0x00,0x01,0x00,0x46,0xff,0xfa,0x04,0x7b,0x04,0x82,0x00,0x1c,0x00,0x00,0x17,0x26,0x35,0x0a,0x01,0x35,0x36,0x37,0x16,0x1f,0x01,0x12,0x25,0x04,0x13,0x14,0x03,0x06,0x23,0x26,0x35,0x12,0x35,0x26,0x27,0x22,0x00,0x03,0x06,0xd8,0x67,0x07,0x24,0x0d,0x58,0x6a,0x07,0x06,0xa8,0x01,0x4f,0x01,0x5d,0x05,0x14,0x0a,0x68,0x55,0x10,0x0a,0x93,0x92,0xfe,0xf4,0x32,0x05,0x02,0x0c,0x68,0x01,0xc3,0x01,0xa2,0x4c,0x5e,0x01,0x09,0x7a,0xf4,0x01,0x6d,0x07,0x0a,0xfe,0x44,0xf2,0xfe,0x98,0x65,0x08,0x63,0x01,0x66,0xdf,0xfd,0x11,0xfe,0x83,0xfe,0x2a,0x5e,0x00,0x00,0x00,0x00,0x02,0x00,0x2d,0xff,0xe9,0x05,0x16,0x04,0x94,0x00,0x0d,0x00,0x19,0x00,0x00,0x01,0x17,0x16,0x00,0x13,0x10,0x00,0x05,0x27,0x24,0x00,0x03,0x36,0x00,0x03,0x12,0x05,0x17,0x24,0x13,0x37,0x34,0x24,0x2f,0x01,0x04,0x02,0x6a,0x4a,0xca,0x01,0x6d,0x2b,0xfe,0xc7,0xfe,0xd7,0x35,0xfe,0xfb,0xfe,0xbc,0x09,0x0e,0x01,0x19,0x5c,0x17,0x01,0x5b,0x51,0x01,0x3b,0x4f,0x0a,0xff,0x00,0xbb,0x33,0xfe,0xc4,0x04,0x94,0x02,0x0d,0xfe,0xe0,0xfe,0xe0,0xfe,0xea,0xfe,0xcd,0x13,0x07,0x1a,0x01,0x41,0x01,0x27,0xe5,0x01,0x2e,0xfd,0xde,0xfe,0xb2,0x61,0x0a,0x1e,0x01,0x0b,0x2f,0xc7,0xee,0x0f,0x01,0x29,0x00,0x00,0x00,0x02,0x00,0x45,0xfd,0xe7,0x04,0xdb,0x04,0x7c,0x00,0x0a,0x00,0x1e,0x00,0x00,0x01,0x06,0x00,0x07,0x17,0x14,0x17,0x36,0x00,0x37,0x26,0x01,0x13,0x06,0x07,0x22,0x27,0x03,0x36,0x37,0x16,0x15,0x17,0x12,0x21,0x04,0x13,0x02,0x00,0x05,0x22,0x03,0x69,0xc0,0xfe,0x94,0x0a,0x03,0xd8,0xad,0x01,0x3f,0x1c,0x06,0xfd,0x2b,0x08,0x0a,0x54,0x67,0x0a,0x2f,0x07,0x5f,0x69,0x06,0xef,0x01,0x75,0x01,0x5a,0x03,0x01,0xfe,0x74,0xfe,0xc4,0x83,0x03,0xbc,0x0c,0xfe,0x8c,0x98,0x56,0x7d,0x0a,0x01,0x01,0x31,0xf0,0xd3,0xfc,0x64,0xfe,0x3b,0x70,0x04,0x77,0x05,0x9d,0x70,0x0a,0x09,0x72,0xef,0x01,0x71,0x12,0xfe,0x81,0xfe,0xf8,0xfe,0x34,0x14,0x00,0x00,0x00,0x02,0x00,0x27,0xfd,0xdd,0x06,0x0a,0x04,0x68,0x00,0x0a,0x00,0x24,0x00,0x00,0x25,0x36,0x00,0x37,0x27,0x34,0x23,0x06,0x00,0x07,0x16,0x00,0x17,0x32,0x36,0x33,0x16,0x17,0x06,0x07,0x24,0x0b,0x01,0x02,0x21,0x24,0x03,0x12,0x00,0x25,0x32,0x17,0x36,0x33,0x32,0x17,0x13,0x01,0x99,0xc0,0x01,0x6c,0x0a,0x03,0xd8,0xad,0xfe,0xc1,0x1c,0x06,0x03,0xd0,0x93,0x22,0x2e,0x19,0x45,0x07,0x01,0xcf,0xfe,0xc4,0x10,0x0b,0xea,0xfe,0x8b,0xfe,0xa6,0x03,0x01,0x01,0x8c,0x01,0x3c,0x96,0x58,0x1e,0x41,0x45,0x13,0x1d,0xaf,0x0c,0x01,0x7e,0x98,0x56,0x7d,0x01,0xfe,0xcf,0xf0,0xd3,0xfd,0xfe,0x01,0x0d,0x0a,0x5a,0x75,0x03,0x28,0x01,0x8a,0x01,0xb3,0xfe,0xad,0x12,0x01,0x7f,0x01,0x08,0x01,0xcc,0x14,0x26,0x26,0x53,0xfb,0x8f,0x00,0x00,0x00,0x01,0x00,0x33,0x00,0x00,0x02,0xfd,0x04,0x89,0x00,0x16,0x00,0x00,0x13,0x16,0x17,0x36,0x37,0x04,0x17,0x06,0x07,0x2e,0x01,0x27,0x06,0x07,0x13,0x06,0x23,0x26,0x27,0x02,0x26,0x35,0x36,0x92,0x63,0x0b,0x41,0x94,0x01,0x12,0x16,0x02,0x47,0x53,0x42,0x43,0xab,0x12,0x1a,0x0e,0x63,0x5a,0x07,0x0c,0x28,0x0e,0x04,0x89,0x06,0x5d,0x53,0x0b,0x12,0xc9,0x59,0x0a,0x01,0x74,0x0a,0x17,0xa0,0xfd,0x6b,0x79,0x01,0x72,0x02,0x99,0xc1,0x5d,0x59,0x00,0x00,0x00,0x00,0x01,0x00,0x45,0xff,0xe9,0x04,0x04,0x04,0x99,0x00,0x20,0x00,0x00,0x01,0x17,0x04,0x17,0x06,0x07,0x2e,0x01,0x23,0x22,0x06,0x07,0x14,0x04,0x13,0x07,0x02,0x05,0x23,0x24,0x27,0x34,0x37,0x32,0x16,0x17,0x24,0x37,0x34,0x24,0x27,0x37,0x12,0x02,0x32,0x45,0x01,0x32,0x0e,0x04,0x46,0x40,0x6d,0x64,0x91,0x9d,0x08,0x02,0xb0,0x2e,0x05,0x38,0xfe,0x5b,0x3a,0xfe,0x70,0x13,0x3c,0x3c,0xa3,0xb8,0x01,0x0b,0x0a,0xfd,0x3e,0x1b,0x02,0x3f,0x04,0x99,0x02,0x15,0xac,0x45,0x0d,0x03,0x4a,0x45,0x54,0x76,0x04,0xfe,0xbe,0x58,0xfe,0xea,0x25,0x1e,0xf5,0x47,0x10,0x8e,0x04,0x07,0x9e,0xad,0x05,0xfc,0x3b,0x01,0x29,0x00,0x00,0x00,0x00,0x01,0x00,0x12,0xff,0xff,0x03,0x78,0x06,0x3e,0x00,0x21,0x00,0x00,0x01,0x16,0x17,0x06,0x2b,0x01,0x27,0x03,0x12,0x17,0x36,0x37,0x36,0x33,0x32,0x15,0x02,0x05,0x24,0x0b,0x01,0x23,0x22,0x27,0x36,0x37,0x33,0x35,0x37,0x36,0x33,0x16,0x17,0x07,0x02,0xd9,0x5a,0x05,0x08,0x5c,0x92,0xbb,0x04,0x02,0xb4,0x69,0x12,0x1d,0x52,0x55,0x2c,0xfe,0xed,0xfe,0x81,0x03,0x01,0x40,0x5c,0x08,0x05,0x5a,0x5d,0x04,0x0c,0x62,0x55,0x0a,0x01,0x05,0x00,0x07,0x5a,0x5b,0x01,0xfd,0x93,0xfe,0xfc,0x09,0x05,0x72,0x5a,0x71,0xfe,0xe3,0x0f,0x0c,0x01,0xd0,0x02,0x69,0x5b,0x5a,0x07,0x01,0xe4,0x59,0x07,0x62,0xd5,0x00,0x00,0x01,0x00,0x35,0x00,0x00,0x04,0x74,0x04,0x8b,0x00,0x1c,0x00,0x00,0x01,0x16,0x15,0x1a,0x01,0x15,0x06,0x07,0x26,0x27,0x03,0x02,0x05,0x24,0x03,0x34,0x13,0x36,0x33,0x16,0x15,0x02,0x15,0x16,0x17,0x32,0x00,0x13,0x36,0x03,0xd8,0x67,0x07,0x2e,0x0d,0x58,0x6a,0x07,0x10,0xa7,0xfe,0xb1,0xfe,0xa3,0x06,0x14,0x0a,0x68,0x55,0x10,0x0a,0x93,0x92,0x01,0x0c,0x32,0x05,0x04,0x87,0x0c,0x68,0xfe,0x3d,0xfe,0x5e,0x4c,0x5e,0x01,0x09,0x7b,0x01,0x07,0xfe,0x79,0x07,0x0a,0x01,0xc2,0xf2,0x01,0x69,0x64,0x08,0x63,0xfe,0x9a,0xdf,0xfd,0x11,0x01,0x7d,0x01,0xd6,0x5e,0x00,0x01,0x00,0x11,0x00,0x04,0x04,0x06,0x04,0x8b,0x00,0x16,0x00,0x00,0x25,0x26,0x27,0x0a,0x01,0x35,0x36,0x37,0x32,0x16,0x13,0x12,0x17,0x36,0x12,0x36,0x33,0x16,0x17,0x14,0x02,0x03,0x06,0x02,0x0f,0x64,0x3f,0xba,0xa1,0x0b,0x54,0x44,0x42,0x70,0x6d,0x3a,0x34,0xe0,0x42,0x4e,0x4a,0x0b,0xa1,0xb9,0x40,0x04,0x01,0xa4,0x01,0xe9,0x01,0x65,0x3a,0x50,0x0a,0x6e,0xfe,0xe4,0xfe,0xea,0x97,0x90,0x02,0x39,0x6e,0x0a,0x50,0x3a,0xfe,0x9b,0xfe,0x17,0xa4,0x00,0x00,0x01,0x00,0x08,0x00,0x04,0x06,0x43,0x04,0x8b,0x00,0x27,0x00,0x00,0x00,0x37,0x16,0x17,0x16,0x12,0x17,0x36,0x12,0x36,0x33,0x16,0x17,0x14,0x02,0x03,0x06,0x07,0x26,0x27,0x02,0x27,0x06,0x03,0x06,0x07,0x26,0x27,0x0a,0x01,0x35,0x36,0x37,0x32,0x16,0x12,0x17,0x36,0x12,0x37,0x02,0xea,0x41,0x36,0x1e,0x21,0xab,0x3a,0x35,0xae,0x42,0x44,0x4a,0x0b,0x89,0x91,0x44,0x5e,0x64,0x3f,0x74,0x4a,0x4b,0x73,0x40,0x5d,0x65,0x43,0x92,0x89,0x0b,0x4a,0x44,0x42,0xab,0x3b,0x34,0xae,0x21,0x04,0x84,0x07,0x07,0x30,0x37,0xfd,0xce,0x97,0x90,0x02,0x39,0x6e,0x0a,0x50,0x3a,0xfe,0x9b,0xfe,0x17,0xa4,0x01,0x01,0xa4,0x01,0xa9,0xbf,0xbf,0xfe,0x57,0xa4,0x01,0x01,0xa4,0x01,0xe9,0x01,0x65,0x3a,0x50,0x0a,0x6e,0xfd,0xce,0x97,0x90,0x02,0x39,0x37,0x00,0x00,0x00,0x01,0x00,0x1c,0x00,0x00,0x04,0x00,0x04,0x80,0x00,0x1f,0x00,0x00,0x09,0x01,0x26,0x27,0x36,0x37,0x16,0x17,0x09,0x01,0x36,0x37,0x16,0x17,0x14,0x07,0x09,0x01,0x16,0x15,0x06,0x07,0x26,0x27,0x09,0x01,0x06,0x07,0x26,0x27,0x36,0x37,0x01,0x8d,0xfe,0xdb,0x4b,0x01,0x06,0x58,0x49,0x32,0x01,0x11,0x01,0x12,0x31,0x4a,0x57,0x06,0x4c,0xfe,0xe3,0x01,0x2d,0x4c,0x06,0x58,0x49,0x31,0xfe,0xe1,0xfe,0xec,0x32,0x49,0x58,0x06,0x01,0x4b,0x02,0x45,0x01,0x4d,0x3b,0x44,0x65,0x0a,0x02,0x56,0xfe,0xd7,0x01,0x29,0x56,0x02,0x0a,0x65,0x44,0x3b,0xfe,0xbc,0xfe,0xa1,0x3a,0x45,0x65,0x0a,0x02,0x57,0x01,0x48,0xfe,0xb7,0x57,0x02,0x0a,0x65,0x45,0x3a,0x00,0x01,0x00,0x32,0xfd,0xe3,0x04,0x55,0x04,0x8b,0x00,0x25,0x00,0x00,0x00,0x05,0x22,0x27,0x26,0x35,0x36,0x37,0x32,0x16,0x33,0x32,0x12,0x11,0x02,0x05,0x24,0x03,0x34,0x13,0x36,0x33,0x16,0x15,0x02,0x15,0x16,0x17,0x32,0x00,0x13,0x36,0x37,0x16,0x15,0x12,0x13,0x10,0x03,0x41,0xfe,0xe3,0x98,0x52,0x3d,0x05,0x3e,0x41,0x51,0x50,0xab,0xbe,0xa8,0xfe,0xb1,0xfe,0xa3,0x05,0x1e,0x0a,0x68,0x55,0x1a,0x0a,0x93,0x92,0x01,0x0c,0x39,0x05,0x66,0x67,0x11,0x01,0xfd,0xe5,0x02,0x29,0x1b,0x4b,0x41,0x1b,0x21,0x01,0x2c,0x01,0xb5,0xfe,0x7f,0x07,0x0a,0x01,0xbc,0xf2,0x01,0x69,0x64,0x08,0x63,0xfe,0x9a,0xdf,0xfd,0x11,0x01,0x7d,0x01,0xd6,0x5e,0x09,0x0c,0x68,0xfe,0x79,0xfe,0xcb,0xfe,0x38,0x00,0x01,0x00,0x32,0x00,0x04,0x03,0x96,0x04,0x7c,0x00,0x15,0x00,0x00,0x01,0x05,0x26,0x27,0x36,0x37,0x21,0x16,0x15,0x14,0x07,0x01,0x21,0x16,0x17,0x06,0x07,0x21,0x26,0x35,0x34,0x37,0x02,0x93,0xfd,0xf5,0x53,0x03,0x0a,0x5f,0x02,0x92,0x69,0x1d,0xfd,0xbc,0x02,0x0b,0x53,0x03,0x0a,0x5f,0xfd,0x6e,0x69,0x1e,0x03,0xb9,0x01,0x11,0x52,0x5b,0x06,0x0f,0x55,0x3a,0x3c,0xfd,0x2a,0x11,0x57,0x57,0x09,0x12,0x55,0x3a,0x3c,0x00,0x00,0x00,0x00,0x01,0x00,0x87,0x02,0xb0,0x03,0x72,0x04,0x0b,0x00,0x17,0x00,0x00,0x00,0x15,0x06,0x07,0x26,0x27,0x26,0x23,0x22,0x07,0x06,0x07,0x26,0x27,0x36,0x37,0x16,0x17,0x16,0x3b,0x01,0x32,0x36,0x37,0x03,0x72,0x2d,0xa6,0x75,0x45,0x48,0x34,0x2b,0x3b,0x15,0x3a,0x2c,0x01,0x2b,0xc3,0x5b,0x49,0x46,0x35,0x04,0x27,0x44,0x3b,0x04,0x02,0x3a,0xca,0x11,0x07,0x19,0x1a,0x4a,0x2c,0x01,0x11,0x3e,0xaa,0x05,0x06,0x19,0x19,0x8e,0x07,0x00,0x00,0xff,0xff,0x00,0x9c,0xfd,0xbd,0x01,0xa0,0x04,0x80,0x00,0x0b,0x00,0x04,0x02,0x6e,0x04,0x7e,0xc0,0x00,0x00,0x02,0x00,0x33,0xff,0xe6,0x04,0x0a,0x07,0x4b,0x00,0x2c,0x00,0x33,0x00,0x00,0x13,0x26,0x03,0x12,0x00,0x25,0x16,0x17,0x13,0x36,0x33,0x16,0x17,0x06,0x07,0x03,0x16,0x17,0x06,0x07,0x26,0x27,0x26,0x27,0x01,0x16,0x17,0x3e,0x02,0x37,0x16,0x17,0x06,0x04,0x07,0x26,0x27,0x07,0x06,0x23,0x26,0x27,0x34,0x37,0x01,0x06,0x07,0x06,0x07,0x16,0x17,0xe2,0xa8,0x07,0x01,0x01,0x1e,0x01,0x14,0x13,0x11,0x9b,0x13,0x3c,0x42,0x01,0x06,0x12,0x78,0xa5,0x03,0x02,0x58,0x35,0x3e,0x12,0x14,0xfe,0xd1,0x26,0x2d,0x8d,0xb8,0x2b,0x47,0x4d,0x06,0x09,0xfe,0xeb,0xdd,0x60,0x4d,0x43,0x1f,0x3a,0x2f,0x06,0x25,0x01,0x87,0x6a,0x62,0x77,0x02,0x09,0x36,0x01,0x20,0x7c,0x01,0x2f,0x01,0x1f,0x01,0x67,0x15,0x01,0x01,0x01,0x8f,0x58,0x05,0x61,0x3c,0x2c,0xfe,0xd3,0x26,0x68,0x53,0x05,0x01,0x1c,0x07,0x06,0xfd,0x0b,0x0c,0x01,0x01,0xa5,0x63,0x01,0x04,0x64,0x74,0xf1,0x05,0x01,0x17,0xa7,0x55,0x04,0x44,0x2c,0x56,0x03,0xee,0x14,0x68,0x80,0xbf,0x94,0x53,0x00,0x00,0x00,0x00,0x01,0x00,0x07,0xff,0xf4,0x05,0xa9,0x07,0x4f,0x00,0x34,0x00,0x00,0x01,0x03,0x05,0x3e,0x01,0x33,0x16,0x17,0x06,0x04,0x07,0x25,0x26,0x27,0x13,0x26,0x27,0x36,0x3f,0x01,0x26,0x27,0x36,0x37,0x12,0x37,0x36,0x25,0x20,0x17,0x16,0x15,0x06,0x23,0x2e,0x01,0x27,0x06,0x07,0x06,0x03,0x21,0x16,0x17,0x06,0x07,0x05,0x07,0x25,0x16,0x17,0x06,0x07,0x01,0x2c,0x28,0x02,0xb3,0xcc,0x89,0x48,0x54,0x01,0x01,0xfe,0xef,0xec,0xfc,0xde,0x53,0x0d,0x2c,0x4c,0x02,0x07,0x56,0x08,0x62,0x03,0x08,0x6d,0x26,0xa8,0xb1,0x01,0x3c,0x01,0x65,0xa1,0x23,0x07,0x57,0x44,0xc9,0xb4,0xc7,0x84,0x77,0x28,0x01,0x50,0x84,0x0c,0x06,0x82,0xfe,0x95,0x07,0x01,0x6a,0x84,0x0c,0x06,0x82,0x02,0xba,0xfe,0x12,0x0c,0x01,0xe9,0x05,0x6a,0x70,0xd6,0x01,0x0b,0x07,0x84,0x02,0x39,0x16,0x49,0x46,0x0e,0x65,0x12,0x53,0x4c,0x09,0x01,0x48,0xb1,0xba,0x07,0x86,0x27,0x3b,0x59,0x07,0x64,0x02,0x01,0x7a,0x61,0xfe,0xf8,0x01,0x58,0x5c,0x0a,0x01,0x5e,0x02,0x02,0x58,0x5b,0x0b,0x00,0x00,0x00,0x02,0x01,0x00,0x05,0x12,0x02,0xde,0x05,0xdc,0x00,0x07,0x00,0x0f,0x00,0x00,0x00,0x15,0x06,0x23,0x22,0x35,0x36,0x37,0x04,0x15,0x06,0x23,0x22,0x35,0x36,0x37,0x01,0xd3,0x14,0x53,0x6c,0x0b,0x52,0x01,0x81,0x13,0x54,0x6c,0x0b,0x52,0x05,0xda,0x6c,0x5c,0x77,0x3f,0x14,0x02,0x6c,0x5c,0x77,0x3f,0x14,0x00,0xff,0xff,0x00,0x16,0x03,0x1e,0x03,0x16,0x07,0x47,0x00,0x63,0x00,0x44,0xff,0xed,0x04,0x88,0x2a,0x3d,0x26,0x66,0x00,0x43,0x00,0x42,0x00,0x5d,0x04,0x41,0x20,0x00,0x40,0x00,0x00,0x00,0x00,0x01,0x00,0x57,0x01,0x13,0x03,0x9f,0x02,0xff,0x00,0x06,0x00,0x00,0x13,0x21,0x11,0x07,0x23,0x11,0x21,0x57,0x03,0x48,0x01,0x62,0xfd,0x1b,0x02,0xff,0xfe,0x15,0x01,0x01,0x88,0x00,0x00,0x01,0x00,0x34,0x05,0x59,0x02,0x9d,0x06,0x0e,0x00,0x0e,0x00,0x00,0x00,0x17,0x06,0x07,0x06,0x0f,0x01,0x26,0x27,0x36,0x33,0x16,0x17,0x36,0x37,0x02,0x93,0x0a,0x05,0x44,0x6d,0x6e,0xd9,0x69,0x03,0x06,0x5d,0x67,0x67,0x65,0x7a,0x06,0x0e,0x4c,0x4d,0x0c,0x0d,0x02,0x01,0x06,0x57,0x4f,0x07,0x01,0x03,0x0e,0x00,0x02,0x00,0x3c,0x03,0x76,0x02,0x68,0x05,0xa2,0x00,0x0b,0x00,0x17,0x00,0x00,0x01,0x22,0x06,0x15,0x14,0x16,0x33,0x32,0x36,0x35,0x34,0x26,0x27,0x32,0x16,0x15,0x14,0x06,0x23,0x22,0x26,0x35,0x34,0x36,0x01,0x53,0x56,0x7b,0x7a,0x57,0x57,0x78,0x79,0x56,0x73,0xa2,0xa4,0x73,0x75,0xa0,0xa3,0x05,0x5c,0x7a,0x57,0x57,0x78,0x78,0x57,0x57,0x7a,0x46,0xa3,0x73,0x72,0xa4,0xa2,0x74,0x74,0xa2,0x00,0x01,0x00,0x28,0xff,0xf6,0x04,0x48,0x05,0xb7,0x00,0x20,0x00,0x00,0x01,0x04,0x13,0x14,0x02,0x05,0x25,0x32,0x16,0x17,0x14,0x23,0x26,0x27,0x04,0x07,0x26,0x35,0x36,0x25,0x24,0x11,0x02,0x25,0x04,0x03,0x06,0x23,0x22,0x27,0x37,0x12,0x25,0x02,0x5c,0x01,0x9b,0x35,0xfa,0xfe,0x7c,0x01,0x0e,0x91,0xf5,0x06,0x6f,0x44,0xd5,0xfe,0x69,0x6f,0x67,0x01,0x01,0x83,0x01,0x9c,0x18,0xfe,0xd9,0xfe,0xf4,0x4c,0x0a,0x5d,0x4c,0x01,0x02,0x44,0x01,0x9a,0x05,0xb7,0x2b,0xfe,0x62,0xe5,0xfe,0xb2,0xe9,0x12,0x30,0x62,0x57,0x19,0x0c,0x11,0x19,0x0a,0x6b,0x6a,0xfc,0xf1,0x01,0x1f,0x01,0x13,0x19,0x0a,0xfe,0xee,0x74,0x6a,0x1f,0x01,0x83,0x2e,0x00,0x00,0x00,0x01,0x00,0x20,0xff,0xf7,0x04,0x57,0x05,0xc5,0x00,0x27,0x00,0x00,0x01,0x04,0x1f,0x01,0x06,0x07,0x04,0x13,0x02,0x05,0x24,0x03,0x36,0x33,0x32,0x12,0x17,0x24,0x37,0x02,0x25,0x06,0x07,0x26,0x35,0x36,0x37,0x36,0x35,0x26,0x27,0x04,0x07,0x14,0x07,0x26,0x27,0x37,0x12,0x25,0x02,0x69,0x01,0x1c,0x3d,0x0a,0x08,0x87,0x01,0x15,0x05,0x33,0xfe,0x16,0xfe,0x00,0x1a,0x0e,0x54,0x42,0x62,0xfb,0x01,0x49,0x23,0x13,0xfe,0xfd,0x5e,0x6c,0x61,0x0b,0xd0,0xcb,0x11,0x86,0xfe,0xbd,0x32,0x5e,0x4c,0x09,0x01,0x49,0x01,0x8f,0x05,0xc5,0x18,0xee,0x3c,0x9e,0x74,0x55,0xfe,0xab,0xfe,0x5d,0x2d,0x04,0x01,0x98,0x47,0xfe,0xfe,0x14,0x0e,0xfb,0x01,0x14,0x0e,0x07,0x07,0x14,0x54,0x5d,0x19,0x18,0xc1,0x72,0x07,0x07,0xc7,0x46,0x0a,0x14,0x55,0x32,0x01,0x20,0x15,0x00,0x00,0x00,0x00,0x01,0x00,0xd3,0x04,0xf2,0x02,0xef,0x06,0x00,0x00,0x0c,0x00,0x00,0x00,0x17,0x14,0x07,0x04,0x23,0x26,0x27,0x34,0x37,0x3e,0x01,0x37,0x02,0xed,0x02,0x54,0xfe,0xab,0x36,0x3c,0x01,0x54,0x9d,0xd9,0x21,0x05,0xf6,0x2c,0x2e,0x1b,0x8f,0x01,0x32,0x31,0x16,0x3b,0x58,0x01,0x00,0x00,0x00,0x00,0x01,0x00,0x9e,0x02,0xa0,0x01,0x7b,0x03,0x83,0x00,0x07,0x00,0x00,0x12,0x37,0x32,0x17,0x14,0x07,0x26,0x27,0x9f,0x64,0x6f,0x09,0x69,0x6c,0x08,0x03,0x7b,0x08,0x6c,0x74,0x03,0x01,0x68,0x00,0x00,0x00,0x00,0x01,0x01,0x58,0xfe,0x3c,0x02,0xe9,0x00,0x08,0x00,0x15,0x00,0x00,0x25,0x33,0x14,0x17,0x16,0x17,0x06,0x07,0x26,0x27,0x36,0x33,0x32,0x16,0x17,0x36,0x37,0x26,0x27,0x26,0x27,0x26,0x01,0xb3,0x6f,0x43,0x82,0x02,0x14,0xac,0xc7,0x0a,0x04,0x31,0x1e,0x29,0x4b,0x50,0x0e,0x07,0x51,0x32,0x27,0x19,0x08,0x67,0x04,0x33,0x80,0x9d,0x11,0x01,0x99,0x2f,0x59,0x08,0x05,0x43,0x4c,0x05,0x0b,0x30,0x21,0x00,0x00,0x00,0x00,0x01,0x00,0xbd,0x00,0x00,0x03,0x27,0x05,0xc1,0x00,0x12,0x00,0x00,0x00,0x17,0x02,0x03,0x06,0x23,0x26,0x27,0x12,0x11,0x06,0x07,0x26,0x27,0x34,0x3f,0x01,0x36,0x33,0x03,0x12,0x15,0x05,0x29,0x09,0x5e,0x57,0x11,0x37,0xe3,0x66,0x48,0x13,0x2f,0xe4,0x8b,0x59,0x05,0xb7,0x40,0xfe,0x08,0xfc,0xc4,0x43,0x03,0x3e,0x03,0x3d,0x01,0x51,0xf9,0x0c,0x07,0x3d,0x48,0x25,0xba,0x8c,0x00,0x00,0x00,0x00,0x04,0x00,0x1b,0xff,0xee,0x06,0x8a,0x05,0xee,0x00,0x12,0x00,0x1d,0x00,0x35,0x00,0x3b,0x00,0x00,0x00,0x17,0x02,0x03,0x06,0x23,0x26,0x27,0x12,0x35,0x06,0x07,0x26,0x27,0x34,0x3f,0x01,0x36,0x33,0x25,0x16,0x17,0x06,0x01,0x26,0x3d,0x01,0x36,0x01,0x36,0x01,0x32,0x17,0x02,0x03,0x37,0x16,0x17,0x06,0x23,0x27,0x17,0x06,0x23,0x26,0x27,0x37,0x06,0x07,0x26,0x3d,0x01,0x36,0x00,0x17,0x00,0x07,0x36,0x37,0x12,0x01,0xa4,0x0e,0x03,0x1b,0x06,0x3e,0x39,0x0c,0x25,0x96,0x43,0x2f,0x0d,0x1f,0x96,0x5c,0x3a,0x02,0x9b,0x36,0x06,0x03,0xfd,0xcc,0x53,0x02,0x02,0x12,0x06,0x01,0xaf,0x44,0x22,0x02,0x18,0x72,0x42,0x0e,0x15,0x25,0x88,0x03,0x0b,0x3b,0x3a,0x07,0x06,0xc5,0xc5,0x45,0x1a,0x01,0xb3,0x1e,0xfe,0xad,0x06,0x93,0xac,0x18,0x05,0xb0,0x2a,0xfe,0xb1,0xfd,0xda,0x2c,0x02,0x29,0x02,0x27,0xdf,0xa5,0x08,0x05,0x28,0x30,0x19,0x7b,0x5d,0x37,0x04,0x65,0x5a,0xfa,0xc3,0x03,0x50,0x21,0x40,0x05,0x06,0x3d,0xfd,0xfc,0x47,0xfe,0xff,0xfe,0xc2,0x07,0x06,0x3e,0x47,0x05,0xa9,0x2b,0x05,0x3d,0x8c,0x01,0x23,0x0a,0x5a,0x1b,0xc7,0x01,0xe9,0x9d,0xfe,0xae,0xb9,0x1e,0x01,0x01,0x49,0x00,0x03,0x00,0x1a,0xff,0xee,0x06,0x40,0x05,0xee,0x00,0x12,0x00,0x1d,0x00,0x3e,0x00,0x00,0x00,0x17,0x02,0x03,0x06,0x23,0x26,0x27,0x12,0x35,0x06,0x07,0x26,0x27,0x34,0x3f,0x01,0x36,0x33,0x25,0x16,0x17,0x06,0x01,0x26,0x3d,0x01,0x36,0x01,0x36,0x01,0x16,0x13,0x14,0x06,0x07,0x37,0x32,0x16,0x17,0x14,0x07,0x26,0x27,0x04,0x07,0x27,0x22,0x27,0x36,0x37,0x24,0x35,0x26,0x27,0x06,0x07,0x14,0x23,0x22,0x27,0x36,0x25,0x01,0xa3,0x0e,0x03,0x1b,0x06,0x3e,0x39,0x0c,0x25,0x96,0x43,0x2f,0x0d,0x1f,0x96,0x5c,0x3a,0x02,0x4c,0x36,0x06,0x03,0xfd,0xcc,0x53,0x02,0x02,0x12,0x06,0x01,0x82,0xff,0x30,0xa3,0xfd,0xb0,0x5e,0xa0,0x04,0x48,0x2d,0x84,0xfe,0xf0,0x3b,0x2b,0x18,0x0d,0x01,0xfc,0x01,0x13,0x1b,0xc0,0xaf,0x47,0x43,0x2a,0x08,0x2e,0x01,0x25,0x05,0xab,0x2a,0xfe,0xb1,0xfd,0xda,0x2c,0x02,0x29,0x02,0x27,0xdf,0xa5,0x08,0x05,0x28,0x30,0x19,0x7b,0x5d,0x3c,0x04,0x65,0x5a,0xfa,0xc3,0x03,0x50,0x21,0x40,0x05,0x06,0x3d,0xfd,0xd7,0x1c,0xfe,0xf3,0x88,0xe6,0x98,0x05,0x18,0x40,0x2c,0x0d,0x11,0x07,0x04,0x17,0x07,0x4c,0x31,0xaa,0x9d,0xbb,0xb3,0x10,0x07,0xab,0x4c,0x52,0xf0,0x31,0x00,0x00,0x00,0x00,0x04,0x00,0x20,0xff,0xd5,0x06,0x8a,0x05,0xd5,0x00,0x27,0x00,0x3f,0x00,0x45,0x00,0x50,0x00,0x00,0x01,0x16,0x1f,0x01,0x06,0x07,0x16,0x17,0x02,0x05,0x24,0x03,0x36,0x33,0x32,0x16,0x17,0x36,0x37,0x26,0x27,0x06,0x07,0x26,0x35,0x36,0x37,0x36,0x35,0x26,0x27,0x06,0x07,0x14,0x07,0x26,0x27,0x35,0x36,0x25,0x01,0x32,0x17,0x02,0x03,0x37,0x16,0x17,0x06,0x23,0x27,0x17,0x06,0x23,0x26,0x27,0x37,0x06,0x07,0x26,0x3d,0x01,0x36,0x00,0x17,0x00,0x07,0x36,0x37,0x12,0x03,0x16,0x17,0x06,0x01,0x26,0x3d,0x01,0x36,0x01,0x36,0x01,0xb4,0xc5,0x2a,0x07,0x06,0x5d,0xc0,0x03,0x23,0xfe,0xad,0xfe,0x9e,0x12,0x18,0x33,0x26,0x44,0xae,0xe3,0x18,0x0d,0xb3,0x41,0x4b,0x43,0x08,0x90,0x8c,0x0c,0x5c,0xe0,0x22,0x41,0x35,0x05,0x32,0x01,0x14,0x04,0x08,0x44,0x22,0x02,0x18,0x72,0x42,0x0e,0x15,0x25,0x88,0x03,0x0b,0x3b,0x3a,0x07,0x06,0xc5,0xc5,0x45,0x1a,0x01,0xb3,0x1e,0xfe,0xad,0x06,0x93,0xac,0x18,0xe4,0x36,0x06,0x03,0xfd,0xcc,0x53,0x02,0x02,0x12,0x06,0x05,0xc5,0x10,0x9c,0x28,0x68,0x4c,0x38,0xe0,0xfe,0xed,0x1e,0x03,0x01,0x0c,0x2f,0xaa,0x0d,0x09,0xa5,0xb5,0x0a,0x05,0x05,0x0e,0x37,0x3d,0x10,0x10,0x7f,0x4b,0x05,0x05,0x83,0x27,0x0d,0x0d,0x31,0x28,0xbd,0x0e,0xfe,0x1d,0x47,0xfe,0xff,0xfe,0xc2,0x07,0x06,0x3e,0x47,0x05,0xa9,0x2b,0x05,0x3d,0x8c,0x01,0x23,0x0a,0x5a,0x1b,0xc7,0x01,0xe9,0x9d,0xfe,0xae,0xb9,0x1e,0x01,0x01,0x49,0x03,0x34,0x04,0x65,0x5a,0xfa,0xc3,0x03,0x50,0x21,0x40,0x05,0x06,0x3d,0x00,0x00,0x00,0x00,0x01,0x00,0x00,0x02,0x1e,0x00,0x01,0x00,0x58,0x01,0x80,0x00,0x06,0x00,0x90,0x00,0x24,0x00,0x37,0xff,0x92,0x00,0x24,0x00,0x3a,0x00,0x6c,0x00,0x24,0x00,0x3c,0xff,0x92,0x00,0x24,0x00,0x59,0x00,0xa0,0x00,0x24,0x00,0x5a,0x00,0xa8,0x00,0x24,0x00,0x5c,0x00,0x5d,0x00,0x29,0x00,0x0f,0xfc,0x7f,0x00,0x29,0x00,0x11,0xfc,0x46,0x00,0x29,0x00,0x24,0x00,0x7e,0x00,0x2f,0x00,0x37,0xfe,0x7e,0x00,0x2f,0x00,0x39,0xfe,0x6a,0x00,0x2f,0x00,0x3a,0xfe,0x66,0x00,0x2f,0x00,0x3c,0xfe,0x47,0x00,0x2f,0x00,0x5c,0x00,0xa3,0x00,0x33,0x00,0x0f,0xfb,0x61,0x00,0x33,0x00,0x11,0xfb,0x28,0x00,0x33,0x00,0x24,0x00,0x62,0x00,0x35,0x00,0x37,0xff,0x3f,0x00,0x35,0x00,0x39,0xff,0xbc,0x00,0x35,0x00,0x3a,0xff,0xbc,0x00,0x35,0x00,0x3c,0xff,0x7d,0x00,0x37,0x00,0x0f,0xfd,0xa3,0x00,0x37,0x00,0x10,0xfe,0x51,0x00,0x37,0x00,0x11,0xfd,0x6a,0x00,0x37,0x00,0x1d,0xfd,0x6a,0x00,0x37,0x00,0x1e,0xfd,0x6a,0x00,0x37,0x00,0x24,0x00,0x36,0x00,0x37,0x00,0x32,0xff,0x28,0x00,0x37,0x00,0x44,0xfd,0xf4,0x00,0x37,0x00,0x46,0xfd,0xdc,0x00,0x37,0x00,0x48,0xfd,0xd5,0x00,0x37,0x00,0x4c,0x00,0x47,0x00,0x37,0x00,0x52,0xfd,0xda,0x00,0x37,0x00,0x55,0xfd,0xd4,0x00,0x37,0x00,0x56,0xfd,0xff,0x00,0x37,0x00,0x58,0xfd,0xe9,0x00,0x37,0x00,0x5a,0xfd,0xdf,0x00,0x37,0x00,0x5c,0xfd,0xdc,0x00,0x39,0x00,0x0f,0xfd,0xd6,0x00,0x39,0x00,0x10,0xff,0x37,0x00,0x39,0x00,0x11,0xfd,0x9d,0x00,0x39,0x00,0x1d,0xff,0x0b,0x00,0x39,0x00,0x1e,0xff,0x0b,0x00,0x39,0x00,0x24,0x00,0x7a,0x00,0x39,0x00,0x44,0xff,0x23,0x00,0x39,0x00,0x48,0xff,0x10,0x00,0x39,0x00,0x4c,0x00,0x34,0x00,0x39,0x00,0x52,0xfe,0xfe,0x00,0x39,0x00,0x55,0xff,0x80,0x00,0x39,0x00,0x58,0xff,0x7d,0x00,0x39,0x00,0x5c,0xff,0x8b,0x00,0x3a,0x00,0x0f,0xfd,0xae,0x00,0x3a,0x00,0x10,0xff,0x34,0x00,0x3a,0x00,0x11,0xfd,0xae,0x00,0x3a,0x00,0x1d,0xff,0x09,0x00,0x3a,0x00,0x1e,0xff,0x09,0x00,0x3a,0x00,0x24,0x00,0x5e,0x00,0x3a,0x00,0x44,0xff,0x13,0x00,0x3a,0x00,0x48,0xff,0x0e,0x00,0x3a,0x00,0x4c,0x00,0x32,0x00,0x3a,0x00,0x52,0xff,0x2f,0x00,0x3a,0x00,0x55,0xff,0x7e,0x00,0x3a,0x00,0x58,0xff,0x7b,0x00,0x3a,0x00,0x5c,0xff,0x89,0x00,0x3c,0x00,0x0f,0xfd,0x95,0x00,0x3c,0x00,0x10,0xfe,0x7e,0x00,0x3c,0x00,0x11,0xfd,0x95,0x00,0x3c,0x00,0x1d,0xfe,0xb1,0x00,0x3c,0x00,0x1e,0xfe,0xb1,0x00,0x3c,0x00,0x24,0x00,0x76,0x00,0x3c,0x00,0x44,0xfe,0x9b,0x00,0x3c,0x00,0x48,0xfe,0x77,0x00,0x3c,0x00,0x4c,0x00,0x56,0x00,0x3c,0x00,0x52,0xfe,0x98,0x00,0x3c,0x00,0x53,0xff,0x1e,0x00,0x3c,0x00,0x54,0xfe,0x40,0x00,0x3c,0x00,0x58,0xff,0x22,0x00,0x3c,0x00,0x59,0xff,0x47,0x00,0x49,0x00,0x48,0xff,0x55,0x00,0x49,0x00,0x49,0x00,0xee,0x00,0x55,0x00,0x0f,0xfe,0x80,0x00,0x55,0x00,0x11,0xfe,0x47,0x00,0x59,0x00,0x0f,0xfe,0x9d,0x00,0x59,0x00,0x11,0xfe,0x64,0x00,0x5a,0x00,0x0f,0xff,0x15,0x00,0x5a,0x00,0x11,0xff,0x21,0x00,0x5c,0x00,0x0f,0xff,0xce,0x00,0x5c,0x00,0x11,0xff,0xce,0x00,0x00,0x00,0x00,0x00,0x2a,0x01,0xfe,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x34,0x00,0x00,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x01,0x00,0x09,0x00,0x3b,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x02,0x00,0x07,0x00,0x34,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x03,0x00,0x16,0x00,0x3b,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x04,0x00,0x09,0x00,0x3b,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x05,0x00,0x2c,0x00,0x51,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x06,0x00,0x08,0x00,0x7d,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x09,0x00,0x0d,0x00,0x85,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x0a,0x00,0x3f,0x00,0x92,0x00,0x01,0x00,0x00,0x00,0x00,0x00,0x0c,0x00,0x19,0x00,0xd1,0x00,0x03,0x00,0x01,0x04,0x03,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x05,0x00,0x02,0x00,0x10,0x00,0xea,0x00,0x03,0x00,0x01,0x04,0x06,0x00,0x02,0x00,0x0c,0x00,0xfa,0x00,0x03,0x00,0x01,0x04,0x07,0x00,0x02,0x00,0x10,0x01,0x06,0x00,0x03,0x00,0x01,0x04,0x08,0x00,0x02,0x00,0x10,0x01,0x16,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x00,0x00,0x96,0x01,0x26,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x01,0x00,0x16,0x01,0x26,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x02,0x00,0x0e,0x01,0xbc,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x03,0x00,0x30,0x01,0xca,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x04,0x00,0x16,0x01,0x26,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x05,0x00,0x6e,0x01,0xfa,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x09,0x00,0x1a,0x01,0x44,0x00,0x03,0x00,0x01,0x04,0x09,0x00,0x0a,0x00,0x7e,0x02,0x68,0x00,0x03,0x00,0x01,0x04,0x0a,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x0b,0x00,0x02,0x00,0x10,0x02,0xe6,0x00,0x03,0x00,0x01,0x04,0x0c,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x0e,0x00,0x02,0x00,0x0c,0x03,0x34,0x00,0x03,0x00,0x01,0x04,0x10,0x00,0x02,0x00,0x0e,0x02,0xf6,0x00,0x03,0x00,0x01,0x04,0x13,0x00,0x02,0x00,0x12,0x03,0x04,0x00,0x03,0x00,0x01,0x04,0x14,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x15,0x00,0x02,0x00,0x10,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x16,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x19,0x00,0x02,0x00,0x0e,0x03,0x26,0x00,0x03,0x00,0x01,0x04,0x1b,0x00,0x02,0x00,0x10,0x03,0x34,0x00,0x03,0x00,0x01,0x04,0x1d,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x1f,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x04,0x24,0x00,0x02,0x00,0x0e,0x03,0x44,0x00,0x03,0x00,0x01,0x04,0x2d,0x00,0x02,0x00,0x0e,0x03,0x52,0x00,0x03,0x00,0x01,0x08,0x0a,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x08,0x16,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x0c,0x0a,0x00,0x02,0x00,0x0c,0x03,0x16,0x00,0x03,0x00,0x01,0x0c,0x0c,0x00,0x02,0x00,0x0c,0x03,0x16,0x54,0x79,0x70,0x65,0x66,0x61,0x63,0x65,0x20,0xa9,0x20,0x28,0x79,0x6f,0x75,0x72,0x20,0x63,0x6f,0x6d,0x70,0x61,0x6e,0x79,0x29,0x2e,0x20,0x32,0x30,0x30,0x38,0x2e,0x20,0x41,0x6c,0x6c,0x20,0x52,0x69,0x67,0x68,0x74,0x73,0x20,0x52,0x65,0x73,0x65,0x72,0x76,0x65,0x64,0x52,0x65,0x67,0x75,0x6c,0x61,0x72,0x51,0x69,0x6b,0x6b,0x69,0x20,0x52,0x65,0x67,0x3a,0x56,0x65,0x72,0x73,0x69,0x6f,0x6e,0x20,0x31,0x2e,0x30,0x30,0x56,0x65,0x72,0x73,0x69,0x6f,0x6e,0x20,0x31,0x2e,0x30,0x30,0x20,0x4d,0x61,0x72,0x63,0x68,0x20,0x32,0x36,0x2c,0x20,0x32,0x30,0x30,0x38,0x2c,0x20,0x69,0x6e,0x69,0x74,0x69,0x61,0x6c,0x20,0x72,0x65,0x6c,0x65,0x61,0x73,0x65,0x51,0x69,0x6b,0x6b,0x69,0x52,0x65,0x67,0x4a,0x6f,0x61,0x6e,0x6e,0x65,0x20,0x54,0x61,0x79,0x6c,0x6f,0x72,0x54,0x68,0x69,0x73,0x20,0x66,0x6f,0x6e,0x74,0x20,0x77,0x61,0x73,0x20,0x63,0x72,0x65,0x61,0x74,0x65,0x64,0x20,0x75,0x73,0x69,0x6e,0x67,0x20,0x46,0x6f,0x6e,0x74,0x43,0x72,0x65,0x61,0x74,0x6f,0x72,0x20,0x35,0x2e,0x36,0x20,0x66,0x72,0x6f,0x6d,0x20,0x48,0x69,0x67,0x68,0x2d,0x4c,0x6f,0x67,0x69,0x63,0x2e,0x63,0x6f,0x6d,0x68,0x74,0x74,0x70,0x3a,0x2f,0x2f,0x77,0x77,0x77,0x2e,0x61,0x72,0x74,0x2d,0x6f,0x66,0x2d,0x71,0x2e,0x63,0x6f,0x2e,0x7a,0x61,0x00,0x6f,0x00,0x62,0x00,0x79,0x01,0x0d,0x00,0x65,0x00,0x6a,0x00,0x6e,0x00,0xe9,0x00,0x6e,0x00,0x6f,0x00,0x72,0x00,0x6d,0x00,0x61,0x00,0x6c,0x00,0x53,0x00,0x74,0x00,0x61,0x00,0x6e,0x00,0x64,0x00,0x61,0x00,0x72,0x00,0x64,0x03,0x9a,0x03,0xb1,0x03,0xbd,0x03,0xbf,0x03,0xbd,0x03,0xb9,0x03,0xba,0x03,0xac,0x00,0x51,0x00,0x61,0x00,0x72,0x00,0x6d,0x00,0x69,0x00,0x63,0x00,0x20,0x00,0x73,0x00,0x61,0x00,0x6e,0x00,0x73,0x00,0x20,0x00,0xa9,0x00,0x20,0x00,0x28,0x00,0x4a,0x00,0x6f,0x00,0x61,0x00,0x6e,0x00,0x6e,0x00,0x65,0x00,0x20,0x00,0x54,0x00,0x61,0x00,0x79,0x00,0x6c,0x00,0x6f,0x00,0x72,0x00,0x20,0x00,0x2d,0x00,0x20,0x00,0x71,0x00,0x61,0x00,0x62,0x00,0x62,0x00,0x6f,0x00,0x6a,0x00,0x6f,0x00,0x40,0x00,0x79,0x00,0x61,0x00,0x68,0x00,0x6f,0x00,0x6f,0x00,0x2e,0x00,0x63,0x00,0x6f,0x00,0x6d,0x00,0x29,0x00,0x20,0x00,0x32,0x00,0x30,0x00,0x30,0x00,0x39,0x00,0x2e,0x00,0x20,0x00,0x41,0x00,0x6c,0x00,0x6c,0x00,0x20,0x00,0x52,0x00,0x69,0x00,0x67,0x00,0x68,0x00,0x74,0x00,0x73,0x00,0x20,0x00,0x52,0x00,0x65,0x00,0x73,0x00,0x65,0x00,0x72,0x00,0x76,0x00,0x65,0x00,0x64,0x00,0x52,0x00,0x65,0x00,0x67,0x00,0x75,0x00,0x6c,0x00,0x61,0x00,0x72,0x00,0x51,0x00,0x61,0x00,0x72,0x00,0x6d,0x00,0x69,0x00,0x63,0x00,0x20,0x00,0x73,0x00,0x61,0x00,0x6e,0x00,0x73,0x00,0x3a,0x00,0x56,0x00,0x65,0x00,0x72,0x00,0x73,0x00,0x69,0x00,0x6f,0x00,0x6e,0x00,0x20,0x00,0x31,0x00,0x2e,0x00,0x30,0x00,0x30,0x00,0x51,0x00,0x61,0x00,0x72,0x00,0x6d,0x00,0x69,0x00,0x63,0x00,0x20,0x00,0x73,0x00,0x61,0x00,0x6e,0x00,0x73,0x00,0x20,0x00,0x56,0x00,0x65,0x00,0x72,0x00,0x73,0x00,0x69,0x00,0x6f,0x00,0x6e,0x00,0x20,0x00,0x31,0x00,0x2e,0x00,0x30,0x00,0x30,0x00,0x3b,0x00,0x20,0x00,0x46,0x00,0x65,0x00,0x62,0x00,0x72,0x00,0x75,0x00,0x61,0x00,0x72,0x00,0x79,0x00,0x20,0x00,0x32,0x00,0x30,0x00,0x30,0x00,0x39,0x00,0x20,0x00,0x69,0x00,0x6e,0x00,0x69,0x00,0x74,0x00,0x69,0x00,0x61,0x00,0x6c,0x00,0x20,0x00,0x72,0x00,0x65,0x00,0x6c,0x00,0x65,0x00,0x61,0x00,0x73,0x00,0x65,0x00,0x54,0x00,0x68,0x00,0x69,0x00,0x73,0x00,0x20,0x00,0x66,0x00,0x6f,0x00,0x6e,0x00,0x74,0x00,0x20,0x00,0x77,0x00,0x61,0x00,0x73,0x00,0x20,0x00,0x63,0x00,0x72,0x00,0x65,0x00,0x61,0x00,0x74,0x00,0x65,0x00,0x64,0x00,0x20,0x00,0x75,0x00,0x73,0x00,0x69,0x00,0x6e,0x00,0x67,0x00,0x20,0x00,0x46,0x00,0x6f,0x00,0x6e,0x00,0x74,0x00,0x43,0x00,0x72,0x00,0x65,0x00,0x61,0x00,0x74,0x00,0x6f,0x00,0x72,0x00,0x20,0x00,0x35,0x00,0x2e,0x00,0x36,0x00,0x20,0x00,0x66,0x00,0x72,0x00,0x6f,0x00,0x6d,0x00,0x20,0x00,0x48,0x00,0x69,0x00,0x67,0x00,0x68,0x00,0x2d,0x00,0x4c,0x00,0x6f,0x00,0x67,0x00,0x69,0x00,0x63,0x00,0x2e,0x00,0x63,0x00,0x6f,0x00,0x6d,0x00,0x4e,0x00,0x6f,0x00,0x72,0x00,0x6d,0x00,0x61,0x00,0x61,0x00,0x6c,0x00,0x69,0x00,0x4e,0x00,0x6f,0x00,0x72,0x00,0x6d,0x00,0x61,0x00,0x6c,0x00,0x65,0x00,0x53,0x00,0x74,0x00,0x61,0x00,0x6e,0x00,0x64,0x00,0x61,0x00,0x61,0x00,0x72,0x00,0x64,0x00,0x4e,0x00,0x6f,0x00,0x72,0x00,0x6d,0x00,0x61,0x00,0x6c,0x00,0x6e,0x00,0x79,0x04,0x1e,0x04,0x31,0x04,0x4b,0x04,0x47,0x04,0x3d,0x04,0x4b,0x04,0x39,0x00,0x4e,0x00,0x6f,0x00,0x72,0x00,0x6d,0x00,0xe1,0x00,0x6c,0x00,0x6e,0x00,0x65,0x00,0x4e,0x00,0x61,0x00,0x76,0x00,0x61,0x00,0x64,0x00,0x6e,0x00,0x6f,0x00,0x41,0x00,0x72,0x00,0x72,0x00,0x75,0x00,0x6e,0x00,0x74,0x00,0x61,0x00,0x00,0x00,0x02,0x00,0x00,0x00,0x00,0x00,0x00,0xff,0x27,0x00,0x96,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x00,0x70,0x00,0x00,0x00,0x01,0x00,0x02,0x00,0x03,0x00,0x04,0x00,0x05,0x00,0x06,0x00,0x07,0x00,0x08,0x00,0x09,0x00,0x0a,0x00,0x0b,0x00,0x0c,0x00,0x0d,0x00,0x0e,0x00,0x0f,0x00,0x10,0x00,0x11,0x00,0x12,0x00,0x13,0x00,0x14,0x00,0x15,0x00,0x16,0x00,0x17,0x00,0x18,0x00,0x19,0x00,0x1a,0x00,0x1b,0x00,0x1c,0x00,0x1d,0x00,0x1e,0x00,0x1f,0x00,0x20,0x00,0x21,0x00,0x22,0x00,0x23,0x00,0x24,0x00,0x25,0x00,0x26,0x00,0x27,0x00,0x28,0x00,0x29,0x00,0x2a,0x00,0x2b,0x00,0x2c,0x00,0x2d,0x00,0x2e,0x00,0x2f,0x00,0x30,0x00,0x31,0x00,0x32,0x00,0x33,0x00,0x34,0x00,0x35,0x00,0x36,0x00,0x37,0x00,0x38,0x00,0x39,0x00,0x3a,0x00,0x3b,0x00,0x3c,0x00,0x3d,0x00,0x3e,0x00,0x3f,0x00,0x40,0x00,0x41,0x00,0x42,0x00,0x43,0x00,0x44,0x00,0x45,0x00,0x46,0x00,0x47,0x00,0x48,0x00,0x49,0x00,0x4a,0x00,0x4b,0x00,0x4c,0x00,0x4d,0x00,0x4e,0x00,0x4f,0x00,0x50,0x00,0x51,0x00,0x52,0x00,0x53,0x00,0x54,0x00,0x55,0x00,0x56,0x00,0x57,0x00,0x58,0x00,0x59,0x00,0x5a,0x00,0x5b,0x00,0x5c,0x00,0x5d,0x00,0x61,0x00,0xa3,0x00,0x84,0x00,0x85,0x00,0x8e,0x00,0x9d,0x00,0xa4,0x00,0xda,0x00,0x83,0x01,0x02,0x01,0x03,0x00,0x8d,0x00,0xc3,0x00,0xde,0x01,0x04,0x00,0xf5,0x00,0xf4,0x00,0xf6,0x07,0x75,0x6e,0x69,0x30,0x30,0x42,0x32,0x07,0x75,0x6e,0x69,0x30,0x30,0x42,0x33,0x07,0x75,0x6e,0x69,0x30,0x30,0x42,0x39,0x00,0x00,0x00,0x00,0x00,0x01,0xff,0xff,0x00,0x02
]
)
