module gx

fn init() {
	eprintln('NB: the `gx` module is deprecated, and will be removed after 2021/12/07.')
	eprintln('All its consts, types, functions are moved into `gg`')
	eprintln('Please `import gg` and replace `gx.` with `gg.` in your source files.')
}
